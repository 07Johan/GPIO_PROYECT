magic
tech sky130A
magscale 1 2
timestamp 1747327185
<< viali >>
rect 5273 20009 5307 20043
rect 8493 20009 8527 20043
rect 9781 20009 9815 20043
rect 11069 20009 11103 20043
rect 11713 20009 11747 20043
rect 13001 20009 13035 20043
rect 14289 20009 14323 20043
rect 17509 20009 17543 20043
rect 17785 20009 17819 20043
rect 10609 19941 10643 19975
rect 18429 19941 18463 19975
rect 5457 19805 5491 19839
rect 5917 19805 5951 19839
rect 6745 19805 6779 19839
rect 7205 19805 7239 19839
rect 8677 19805 8711 19839
rect 9167 19805 9201 19839
rect 9321 19805 9355 19839
rect 9965 19805 9999 19839
rect 10425 19805 10459 19839
rect 10885 19805 10919 19839
rect 11253 19805 11287 19839
rect 11897 19805 11931 19839
rect 13185 19805 13219 19839
rect 13829 19805 13863 19839
rect 14473 19805 14507 19839
rect 14933 19805 14967 19839
rect 16221 19805 16255 19839
rect 17325 19805 17359 19839
rect 17601 19805 17635 19839
rect 17877 19805 17911 19839
rect 18337 19805 18371 19839
rect 18613 19805 18647 19839
rect 6101 19669 6135 19703
rect 6561 19669 6595 19703
rect 7389 19669 7423 19703
rect 8953 19669 8987 19703
rect 10701 19669 10735 19703
rect 13645 19669 13679 19703
rect 15117 19669 15151 19703
rect 16405 19669 16439 19703
rect 18061 19669 18095 19703
rect 18153 19669 18187 19703
rect 4445 19465 4479 19499
rect 4905 19465 4939 19499
rect 6561 19465 6595 19499
rect 9505 19465 9539 19499
rect 11345 19465 11379 19499
rect 11713 19465 11747 19499
rect 13277 19465 13311 19499
rect 13829 19465 13863 19499
rect 14933 19465 14967 19499
rect 18521 19465 18555 19499
rect 2697 19329 2731 19363
rect 4721 19329 4755 19363
rect 5641 19329 5675 19363
rect 5733 19329 5767 19363
rect 5917 19329 5951 19363
rect 7205 19329 7239 19363
rect 7757 19329 7791 19363
rect 9597 19329 9631 19363
rect 11529 19329 11563 19363
rect 12908 19329 12942 19363
rect 13001 19329 13035 19363
rect 13093 19329 13127 19363
rect 13645 19329 13679 19363
rect 15209 19329 15243 19363
rect 15393 19329 15427 19363
rect 18705 19329 18739 19363
rect 2973 19261 3007 19295
rect 8033 19261 8067 19295
rect 9873 19261 9907 19295
rect 16681 19261 16715 19295
rect 16957 19261 16991 19295
rect 6929 19193 6963 19227
rect 14565 19193 14599 19227
rect 15117 19193 15151 19227
rect 5549 19125 5583 19159
rect 5825 19125 5859 19159
rect 6377 19125 6411 19159
rect 6561 19125 6595 19159
rect 7297 19125 7331 19159
rect 12817 19125 12851 19159
rect 14933 19125 14967 19159
rect 15301 19125 15335 19159
rect 18429 19125 18463 19159
rect 3893 18921 3927 18955
rect 8217 18921 8251 18955
rect 8953 18921 8987 18955
rect 9781 18921 9815 18955
rect 10517 18921 10551 18955
rect 10701 18921 10735 18955
rect 11621 18921 11655 18955
rect 13737 18921 13771 18955
rect 16957 18921 16991 18955
rect 18061 18921 18095 18955
rect 10149 18853 10183 18887
rect 18153 18853 18187 18887
rect 4353 18785 4387 18819
rect 6193 18785 6227 18819
rect 7941 18785 7975 18819
rect 11989 18785 12023 18819
rect 14105 18785 14139 18819
rect 1409 18717 1443 18751
rect 1777 18717 1811 18751
rect 3985 18717 4019 18751
rect 8033 18717 8067 18751
rect 9229 18717 9263 18751
rect 9321 18717 9355 18751
rect 9413 18717 9447 18751
rect 9597 18717 9631 18751
rect 9873 18717 9907 18751
rect 11713 18717 11747 18751
rect 16619 18717 16653 18751
rect 16773 18717 16807 18751
rect 16865 18717 16899 18751
rect 17877 18717 17911 18751
rect 18337 18717 18371 18751
rect 18429 18717 18463 18751
rect 2053 18649 2087 18683
rect 4629 18649 4663 18683
rect 6469 18649 6503 18683
rect 10517 18649 10551 18683
rect 12265 18649 12299 18683
rect 14381 18649 14415 18683
rect 1593 18581 1627 18615
rect 3525 18581 3559 18615
rect 6101 18581 6135 18615
rect 15853 18581 15887 18615
rect 16405 18581 16439 18615
rect 18613 18581 18647 18615
rect 1593 18377 1627 18411
rect 1777 18377 1811 18411
rect 2329 18377 2363 18411
rect 2697 18377 2731 18411
rect 2881 18377 2915 18411
rect 3249 18377 3283 18411
rect 5549 18377 5583 18411
rect 5917 18377 5951 18411
rect 9413 18377 9447 18411
rect 12173 18377 12207 18411
rect 13093 18377 13127 18411
rect 14657 18377 14691 18411
rect 15025 18377 15059 18411
rect 18429 18377 18463 18411
rect 18797 18377 18831 18411
rect 7205 18309 7239 18343
rect 2513 18241 2547 18275
rect 2789 18241 2823 18275
rect 2881 18241 2915 18275
rect 3065 18241 3099 18275
rect 3341 18241 3375 18275
rect 5733 18241 5767 18275
rect 6009 18241 6043 18275
rect 6561 18241 6595 18275
rect 7297 18241 7331 18275
rect 7481 18241 7515 18275
rect 7573 18241 7607 18275
rect 7665 18241 7699 18275
rect 8247 18241 8281 18275
rect 8401 18241 8435 18275
rect 9229 18241 9263 18275
rect 12403 18241 12437 18275
rect 12538 18247 12572 18281
rect 12633 18244 12667 18278
rect 12817 18241 12851 18275
rect 13001 18241 13035 18275
rect 14841 18241 14875 18275
rect 15117 18241 15151 18275
rect 15393 18241 15427 18275
rect 15577 18241 15611 18275
rect 18613 18241 18647 18275
rect 6745 18173 6779 18207
rect 8033 18173 8067 18207
rect 15761 18173 15795 18207
rect 16681 18173 16715 18207
rect 16957 18173 16991 18207
rect 2145 18105 2179 18139
rect 15301 18105 15335 18139
rect 1777 18037 1811 18071
rect 7941 18037 7975 18071
rect 16221 18037 16255 18071
rect 1593 17833 1627 17867
rect 12357 17833 12391 17867
rect 16957 17833 16991 17867
rect 17693 17833 17727 17867
rect 6745 17765 6779 17799
rect 11805 17697 11839 17731
rect 15577 17697 15611 17731
rect 1409 17629 1443 17663
rect 6377 17629 6411 17663
rect 6470 17629 6504 17663
rect 8585 17629 8619 17663
rect 10609 17629 10643 17663
rect 10885 17629 10919 17663
rect 11161 17629 11195 17663
rect 11989 17629 12023 17663
rect 15853 17629 15887 17663
rect 16313 17629 16347 17663
rect 16497 17629 16531 17663
rect 16589 17629 16623 17663
rect 16681 17629 16715 17663
rect 17601 17629 17635 17663
rect 18797 17629 18831 17663
rect 8677 17493 8711 17527
rect 10425 17493 10459 17527
rect 10793 17493 10827 17527
rect 11069 17493 11103 17527
rect 14105 17493 14139 17527
rect 18613 17493 18647 17527
rect 9321 17289 9355 17323
rect 11529 17289 11563 17323
rect 11897 17289 11931 17323
rect 14749 17289 14783 17323
rect 15485 17289 15519 17323
rect 3433 17221 3467 17255
rect 6561 17221 6595 17255
rect 7849 17221 7883 17255
rect 9873 17221 9907 17255
rect 1593 17153 1627 17187
rect 2329 17153 2363 17187
rect 2421 17153 2455 17187
rect 2513 17153 2547 17187
rect 2697 17153 2731 17187
rect 4077 17153 4111 17187
rect 6193 17153 6227 17187
rect 7573 17153 7607 17187
rect 9597 17153 9631 17187
rect 11529 17153 11563 17187
rect 11713 17153 11747 17187
rect 12172 17153 12206 17187
rect 12265 17153 12299 17187
rect 14841 17153 14875 17187
rect 15117 17153 15151 17187
rect 15210 17153 15244 17187
rect 17509 17153 17543 17187
rect 17601 17153 17635 17187
rect 17693 17153 17727 17187
rect 17877 17153 17911 17187
rect 18183 17153 18217 17187
rect 18337 17153 18371 17187
rect 18429 17153 18463 17187
rect 3893 17085 3927 17119
rect 11345 17085 11379 17119
rect 17969 17085 18003 17119
rect 1409 16949 1443 16983
rect 2053 16949 2087 16983
rect 6101 16949 6135 16983
rect 17233 16949 17267 16983
rect 18521 16949 18555 16983
rect 1409 16745 1443 16779
rect 6469 16745 6503 16779
rect 18797 16745 18831 16779
rect 4261 16677 4295 16711
rect 1685 16609 1719 16643
rect 1961 16609 1995 16643
rect 4721 16609 4755 16643
rect 4997 16609 5031 16643
rect 6561 16609 6595 16643
rect 10701 16609 10735 16643
rect 10977 16609 11011 16643
rect 17049 16609 17083 16643
rect 17325 16609 17359 16643
rect 1593 16541 1627 16575
rect 3985 16541 4019 16575
rect 4536 16541 4570 16575
rect 4629 16541 4663 16575
rect 8953 16541 8987 16575
rect 9107 16541 9141 16575
rect 12725 16541 12759 16575
rect 14105 16541 14139 16575
rect 14289 16541 14323 16575
rect 14473 16541 14507 16575
rect 14933 16541 14967 16575
rect 15026 16541 15060 16575
rect 8309 16473 8343 16507
rect 12633 16473 12667 16507
rect 3433 16405 3467 16439
rect 4077 16405 4111 16439
rect 9321 16405 9355 16439
rect 12449 16405 12483 16439
rect 14197 16405 14231 16439
rect 14565 16405 14599 16439
rect 15301 16405 15335 16439
rect 2421 16201 2455 16235
rect 2789 16201 2823 16235
rect 4905 16201 4939 16235
rect 9229 16201 9263 16235
rect 15485 16201 15519 16235
rect 18429 16201 18463 16235
rect 7757 16133 7791 16167
rect 1409 16065 1443 16099
rect 2053 16065 2087 16099
rect 2146 16065 2180 16099
rect 2697 16065 2731 16099
rect 3157 16065 3191 16099
rect 7205 16065 7239 16099
rect 7389 16065 7423 16099
rect 9505 16065 9539 16099
rect 14197 16065 14231 16099
rect 16681 16065 16715 16099
rect 18797 16065 18831 16099
rect 3433 15997 3467 16031
rect 7481 15997 7515 16031
rect 9321 15997 9355 16031
rect 12357 15997 12391 16031
rect 12633 15997 12667 16031
rect 16957 15997 16991 16031
rect 9689 15929 9723 15963
rect 1593 15861 1627 15895
rect 7297 15861 7331 15895
rect 14105 15861 14139 15895
rect 18613 15861 18647 15895
rect 8033 15657 8067 15691
rect 8585 15657 8619 15691
rect 10793 15657 10827 15691
rect 13369 15657 13403 15691
rect 14197 15657 14231 15691
rect 17141 15657 17175 15691
rect 17509 15657 17543 15691
rect 2329 15589 2363 15623
rect 16681 15589 16715 15623
rect 6285 15521 6319 15555
rect 9045 15521 9079 15555
rect 15669 15521 15703 15555
rect 15945 15521 15979 15555
rect 16221 15521 16255 15555
rect 1593 15453 1627 15487
rect 2513 15453 2547 15487
rect 5825 15453 5859 15487
rect 8309 15453 8343 15487
rect 8493 15453 8527 15487
rect 11069 15453 11103 15487
rect 13001 15453 13035 15487
rect 13277 15453 13311 15487
rect 16037 15453 16071 15487
rect 16773 15453 16807 15487
rect 17417 15453 17451 15487
rect 18613 15453 18647 15487
rect 6561 15385 6595 15419
rect 8217 15385 8251 15419
rect 9321 15385 9355 15419
rect 10977 15385 11011 15419
rect 17141 15385 17175 15419
rect 1409 15317 1443 15351
rect 5733 15317 5767 15351
rect 17325 15317 17359 15351
rect 18797 15317 18831 15351
rect 3157 15113 3191 15147
rect 7113 15113 7147 15147
rect 7205 15113 7239 15147
rect 7573 15113 7607 15147
rect 14105 15113 14139 15147
rect 14473 15113 14507 15147
rect 6929 15045 6963 15079
rect 11713 15045 11747 15079
rect 1409 14977 1443 15011
rect 3525 14977 3559 15011
rect 3709 14977 3743 15011
rect 3801 14977 3835 15011
rect 5641 14977 5675 15011
rect 7389 14977 7423 15011
rect 7665 14977 7699 15011
rect 11805 14977 11839 15011
rect 14289 14977 14323 15011
rect 14565 14977 14599 15011
rect 17417 14977 17451 15011
rect 17509 14977 17543 15011
rect 17601 14977 17635 15011
rect 17785 14977 17819 15011
rect 18152 14977 18186 15011
rect 18245 14977 18279 15011
rect 18797 14977 18831 15011
rect 1685 14909 1719 14943
rect 4077 14909 4111 14943
rect 6561 14909 6595 14943
rect 15485 14909 15519 14943
rect 15669 14909 15703 14943
rect 16129 14909 16163 14943
rect 17877 14909 17911 14943
rect 3617 14773 3651 14807
rect 5549 14773 5583 14807
rect 6929 14773 6963 14807
rect 17141 14773 17175 14807
rect 18613 14773 18647 14807
rect 2513 14569 2547 14603
rect 3801 14569 3835 14603
rect 2237 14501 2271 14535
rect 4353 14501 4387 14535
rect 1501 14433 1535 14467
rect 5089 14433 5123 14467
rect 14756 14433 14790 14467
rect 15025 14433 15059 14467
rect 17325 14433 17359 14467
rect 1777 14365 1811 14399
rect 2421 14365 2455 14399
rect 3985 14365 4019 14399
rect 4261 14365 4295 14399
rect 4353 14365 4387 14399
rect 4537 14365 4571 14399
rect 6837 14365 6871 14399
rect 14289 14365 14323 14399
rect 14473 14365 14507 14399
rect 14657 14365 14691 14399
rect 17049 14365 17083 14399
rect 2237 14297 2271 14331
rect 4169 14297 4203 14331
rect 1685 14229 1719 14263
rect 14197 14229 14231 14263
rect 14473 14229 14507 14263
rect 16497 14229 16531 14263
rect 18797 14229 18831 14263
rect 1777 14025 1811 14059
rect 17049 14025 17083 14059
rect 18061 14025 18095 14059
rect 18797 14025 18831 14059
rect 5365 13957 5399 13991
rect 5641 13957 5675 13991
rect 1501 13889 1535 13923
rect 1961 13889 1995 13923
rect 3157 13889 3191 13923
rect 3525 13889 3559 13923
rect 4169 13889 4203 13923
rect 4353 13889 4387 13923
rect 4997 13889 5031 13923
rect 5151 13889 5185 13923
rect 13369 13889 13403 13923
rect 16681 13889 16715 13923
rect 17969 13889 18003 13923
rect 18613 13889 18647 13923
rect 3617 13821 3651 13855
rect 5549 13821 5583 13855
rect 5825 13821 5859 13855
rect 1685 13753 1719 13787
rect 3065 13685 3099 13719
rect 4353 13685 4387 13719
rect 17049 13685 17083 13719
rect 17233 13685 17267 13719
rect 3801 13481 3835 13515
rect 6101 13481 6135 13515
rect 15393 13481 15427 13515
rect 16037 13481 16071 13515
rect 18613 13481 18647 13515
rect 1869 13345 1903 13379
rect 4353 13345 4387 13379
rect 4629 13345 4663 13379
rect 16589 13345 16623 13379
rect 18061 13345 18095 13379
rect 1777 13277 1811 13311
rect 4077 13277 4111 13311
rect 4261 13277 4295 13311
rect 6377 13277 6411 13311
rect 13645 13277 13679 13311
rect 13829 13277 13863 13311
rect 13921 13277 13955 13311
rect 14105 13277 14139 13311
rect 16129 13277 16163 13311
rect 16313 13277 16347 13311
rect 18337 13277 18371 13311
rect 18429 13277 18463 13311
rect 2145 13209 2179 13243
rect 6285 13209 6319 13243
rect 18245 13209 18279 13243
rect 1593 13141 1627 13175
rect 3617 13141 3651 13175
rect 3985 13141 4019 13175
rect 13461 13141 13495 13175
rect 1409 12937 1443 12971
rect 2605 12937 2639 12971
rect 14657 12937 14691 12971
rect 15669 12937 15703 12971
rect 18337 12937 18371 12971
rect 18613 12937 18647 12971
rect 1593 12801 1627 12835
rect 1685 12801 1719 12835
rect 2789 12801 2823 12835
rect 2881 12801 2915 12835
rect 3065 12801 3099 12835
rect 3249 12801 3283 12835
rect 12909 12801 12943 12835
rect 15301 12801 15335 12835
rect 15455 12801 15489 12835
rect 18153 12801 18187 12835
rect 18797 12801 18831 12835
rect 2973 12733 3007 12767
rect 13185 12733 13219 12767
rect 1869 12597 1903 12631
rect 13921 12257 13955 12291
rect 14105 12257 14139 12291
rect 18060 12189 18094 12223
rect 18153 12189 18187 12223
rect 18797 12189 18831 12223
rect 11897 12121 11931 12155
rect 13645 12121 13679 12155
rect 14381 12121 14415 12155
rect 15853 12053 15887 12087
rect 17785 12053 17819 12087
rect 18613 12053 18647 12087
rect 13001 11849 13035 11883
rect 15117 11849 15151 11883
rect 18705 11849 18739 11883
rect 1685 11781 1719 11815
rect 9321 11781 9355 11815
rect 16497 11781 16531 11815
rect 3985 11713 4019 11747
rect 4077 11713 4111 11747
rect 4169 11713 4203 11747
rect 4353 11713 4387 11747
rect 4445 11713 4479 11747
rect 4813 11713 4847 11747
rect 4997 11713 5031 11747
rect 5457 11713 5491 11747
rect 13093 11713 13127 11747
rect 15025 11713 15059 11747
rect 15393 11713 15427 11747
rect 15547 11713 15581 11747
rect 15761 11713 15795 11747
rect 16037 11713 16071 11747
rect 16957 11713 16991 11747
rect 1409 11645 1443 11679
rect 4721 11645 4755 11679
rect 15853 11645 15887 11679
rect 17233 11645 17267 11679
rect 3157 11509 3191 11543
rect 3709 11509 3743 11543
rect 4537 11509 4571 11543
rect 4905 11509 4939 11543
rect 5089 11509 5123 11543
rect 5365 11509 5399 11543
rect 10609 11509 10643 11543
rect 2145 11305 2179 11339
rect 3249 11305 3283 11339
rect 4353 11305 4387 11339
rect 5181 11305 5215 11339
rect 5273 11305 5307 11339
rect 16589 11305 16623 11339
rect 17141 11305 17175 11339
rect 18061 11305 18095 11339
rect 3157 11237 3191 11271
rect 16221 11237 16255 11271
rect 3525 11169 3559 11203
rect 4721 11169 4755 11203
rect 4997 11169 5031 11203
rect 5181 11169 5215 11203
rect 5549 11169 5583 11203
rect 7297 11169 7331 11203
rect 1409 11101 1443 11135
rect 2237 11101 2271 11135
rect 3617 11101 3651 11135
rect 3893 11101 3927 11135
rect 4169 11101 4203 11135
rect 4445 11101 4479 11135
rect 4905 11101 4939 11135
rect 5365 11101 5399 11135
rect 7573 11101 7607 11135
rect 15301 11101 15335 11135
rect 15485 11101 15519 11135
rect 15761 11101 15795 11135
rect 17417 11101 17451 11135
rect 17509 11101 17543 11135
rect 17601 11101 17635 11135
rect 17785 11101 17819 11135
rect 17969 11101 18003 11135
rect 18797 11101 18831 11135
rect 2789 11033 2823 11067
rect 4537 11033 4571 11067
rect 5825 11033 5859 11067
rect 7481 11033 7515 11067
rect 15669 11033 15703 11067
rect 16589 11033 16623 11067
rect 1593 10965 1627 10999
rect 3985 10965 4019 10999
rect 15485 10965 15519 10999
rect 16773 10965 16807 10999
rect 18613 10965 18647 10999
rect 3157 10761 3191 10795
rect 6377 10761 6411 10795
rect 6837 10761 6871 10795
rect 16037 10761 16071 10795
rect 1685 10693 1719 10727
rect 5549 10693 5583 10727
rect 6745 10693 6779 10727
rect 5825 10625 5859 10659
rect 18153 10625 18187 10659
rect 18613 10625 18647 10659
rect 1409 10557 1443 10591
rect 4077 10557 4111 10591
rect 6929 10557 6963 10591
rect 14289 10557 14323 10591
rect 14565 10557 14599 10591
rect 18337 10421 18371 10455
rect 18797 10421 18831 10455
rect 2421 10217 2455 10251
rect 15209 10217 15243 10251
rect 18337 10217 18371 10251
rect 1409 10081 1443 10115
rect 1685 10081 1719 10115
rect 16865 10081 16899 10115
rect 2329 10013 2363 10047
rect 15393 10013 15427 10047
rect 15577 10013 15611 10047
rect 15669 10013 15703 10047
rect 16589 10013 16623 10047
rect 18429 10013 18463 10047
rect 18521 9945 18555 9979
rect 1593 9673 1627 9707
rect 2145 9605 2179 9639
rect 4169 9605 4203 9639
rect 5825 9605 5859 9639
rect 13185 9605 13219 9639
rect 1409 9537 1443 9571
rect 1869 9537 1903 9571
rect 5917 9537 5951 9571
rect 11989 9537 12023 9571
rect 18705 9537 18739 9571
rect 3893 9469 3927 9503
rect 16681 9469 16715 9503
rect 16957 9469 16991 9503
rect 18429 9469 18463 9503
rect 12173 9401 12207 9435
rect 3617 9333 3651 9367
rect 5641 9333 5675 9367
rect 14473 9333 14507 9367
rect 18521 9333 18555 9367
rect 2973 9129 3007 9163
rect 17325 9129 17359 9163
rect 18797 9129 18831 9163
rect 1409 9061 1443 9095
rect 9597 8993 9631 9027
rect 9965 8993 9999 9027
rect 1593 8925 1627 8959
rect 1961 8925 1995 8959
rect 2881 8925 2915 8959
rect 5733 8925 5767 8959
rect 8953 8925 8987 8959
rect 9137 8925 9171 8959
rect 9229 8925 9263 8959
rect 9321 8925 9355 8959
rect 9689 8925 9723 8959
rect 11713 8925 11747 8959
rect 14197 8925 14231 8959
rect 16221 8925 16255 8959
rect 17233 8925 17267 8959
rect 18337 8925 18371 8959
rect 18613 8925 18647 8959
rect 11621 8857 11655 8891
rect 14473 8857 14507 8891
rect 16129 8857 16163 8891
rect 1777 8789 1811 8823
rect 11437 8789 11471 8823
rect 15945 8789 15979 8823
rect 18521 8789 18555 8823
rect 4169 8585 4203 8619
rect 4537 8585 4571 8619
rect 9413 8585 9447 8619
rect 6377 8517 6411 8551
rect 16221 8517 16255 8551
rect 3157 8449 3191 8483
rect 4261 8449 4295 8483
rect 4629 8449 4663 8483
rect 8125 8449 8159 8483
rect 9627 8449 9661 8483
rect 9781 8449 9815 8483
rect 13185 8449 13219 8483
rect 16865 8449 16899 8483
rect 2881 8381 2915 8415
rect 3801 8381 3835 8415
rect 15577 8381 15611 8415
rect 15761 8381 15795 8415
rect 17141 8381 17175 8415
rect 3985 8313 4019 8347
rect 1409 8245 1443 8279
rect 18613 8245 18647 8279
rect 1409 8041 1443 8075
rect 2329 8041 2363 8075
rect 16129 8041 16163 8075
rect 17049 8041 17083 8075
rect 18337 8041 18371 8075
rect 4169 7973 4203 8007
rect 3893 7905 3927 7939
rect 3985 7905 4019 7939
rect 4261 7905 4295 7939
rect 14105 7905 14139 7939
rect 1593 7837 1627 7871
rect 1685 7837 1719 7871
rect 2053 7837 2087 7871
rect 2421 7837 2455 7871
rect 2697 7837 2731 7871
rect 3801 7837 3835 7871
rect 9137 7837 9171 7871
rect 13737 7837 13771 7871
rect 15945 7837 15979 7871
rect 16038 7837 16072 7871
rect 17325 7837 17359 7871
rect 17417 7837 17451 7871
rect 17509 7837 17543 7871
rect 17693 7837 17727 7871
rect 18060 7837 18094 7871
rect 18153 7837 18187 7871
rect 18429 7837 18463 7871
rect 18613 7837 18647 7871
rect 1869 7769 1903 7803
rect 4099 7769 4133 7803
rect 4537 7769 4571 7803
rect 14381 7769 14415 7803
rect 17785 7769 17819 7803
rect 2513 7701 2547 7735
rect 6009 7701 6043 7735
rect 9045 7701 9079 7735
rect 13829 7701 13863 7735
rect 15853 7701 15887 7735
rect 18797 7701 18831 7735
rect 1409 7497 1443 7531
rect 3341 7497 3375 7531
rect 4721 7497 4755 7531
rect 5457 7497 5491 7531
rect 14657 7497 14691 7531
rect 15025 7497 15059 7531
rect 15209 7497 15243 7531
rect 4445 7429 4479 7463
rect 8033 7429 8067 7463
rect 15853 7429 15887 7463
rect 1593 7361 1627 7395
rect 3617 7361 3651 7395
rect 3709 7361 3743 7395
rect 3801 7361 3835 7395
rect 3985 7361 4019 7395
rect 4261 7361 4295 7395
rect 4537 7361 4571 7395
rect 4813 7361 4847 7395
rect 5549 7361 5583 7395
rect 6745 7361 6779 7395
rect 6837 7361 6871 7395
rect 7389 7361 7423 7395
rect 12909 7361 12943 7395
rect 14841 7361 14875 7395
rect 15117 7361 15151 7395
rect 15209 7361 15243 7395
rect 15393 7361 15427 7395
rect 15485 7361 15519 7395
rect 18153 7361 18187 7395
rect 18613 7361 18647 7395
rect 6929 7293 6963 7327
rect 7757 7293 7791 7327
rect 9597 7293 9631 7327
rect 9781 7293 9815 7327
rect 16037 7225 16071 7259
rect 4077 7157 4111 7191
rect 6377 7157 6411 7191
rect 7297 7157 7331 7191
rect 9505 7157 9539 7191
rect 9965 7157 9999 7191
rect 15853 7157 15887 7191
rect 18337 7157 18371 7191
rect 18797 7157 18831 7191
rect 3985 6953 4019 6987
rect 5812 6953 5846 6987
rect 7297 6953 7331 6987
rect 12436 6953 12470 6987
rect 14105 6953 14139 6987
rect 15840 6953 15874 6987
rect 18337 6953 18371 6987
rect 18613 6953 18647 6987
rect 9413 6885 9447 6919
rect 4077 6817 4111 6851
rect 5549 6817 5583 6851
rect 12173 6817 12207 6851
rect 14749 6817 14783 6851
rect 17325 6817 17359 6851
rect 1409 6749 1443 6783
rect 3801 6749 3835 6783
rect 3893 6749 3927 6783
rect 4169 6749 4203 6783
rect 8401 6749 8435 6783
rect 8585 6749 8619 6783
rect 9045 6749 9079 6783
rect 9199 6749 9233 6783
rect 14289 6749 14323 6783
rect 14565 6749 14599 6783
rect 14841 6749 14875 6783
rect 15577 6749 15611 6783
rect 18153 6749 18187 6783
rect 18429 6749 18463 6783
rect 1685 6681 1719 6715
rect 3157 6613 3191 6647
rect 8585 6613 8619 6647
rect 13921 6613 13955 6647
rect 14473 6613 14507 6647
rect 2421 6409 2455 6443
rect 3433 6409 3467 6443
rect 9321 6409 9355 6443
rect 14473 6409 14507 6443
rect 16773 6409 16807 6443
rect 18613 6409 18647 6443
rect 9505 6341 9539 6375
rect 12541 6341 12575 6375
rect 1501 6273 1535 6307
rect 1777 6273 1811 6307
rect 2329 6273 2363 6307
rect 2973 6273 3007 6307
rect 9597 6273 9631 6307
rect 14381 6273 14415 6307
rect 14565 6273 14599 6307
rect 14841 6273 14875 6307
rect 16865 6273 16899 6307
rect 17968 6273 18002 6307
rect 18061 6273 18095 6307
rect 18797 6273 18831 6307
rect 7573 6205 7607 6239
rect 7849 6205 7883 6239
rect 15025 6205 15059 6239
rect 1685 6137 1719 6171
rect 3341 6137 3375 6171
rect 17693 6137 17727 6171
rect 1961 6069 1995 6103
rect 13829 6069 13863 6103
rect 15485 6069 15519 6103
rect 8401 5865 8435 5899
rect 8953 5865 8987 5899
rect 15589 5865 15623 5899
rect 16405 5865 16439 5899
rect 16589 5865 16623 5899
rect 18613 5865 18647 5899
rect 2237 5797 2271 5831
rect 8217 5797 8251 5831
rect 16037 5797 16071 5831
rect 4077 5729 4111 5763
rect 15853 5729 15887 5763
rect 16865 5729 16899 5763
rect 1593 5661 1627 5695
rect 1869 5661 1903 5695
rect 2145 5661 2179 5695
rect 2329 5661 2363 5695
rect 2421 5661 2455 5695
rect 2605 5661 2639 5695
rect 3801 5661 3835 5695
rect 3985 5661 4019 5695
rect 6101 5661 6135 5695
rect 8125 5661 8159 5695
rect 8769 5661 8803 5695
rect 9137 5661 9171 5695
rect 9321 5661 9355 5695
rect 9413 5661 9447 5695
rect 11069 5661 11103 5695
rect 12356 5661 12390 5695
rect 12449 5661 12483 5695
rect 12541 5661 12575 5695
rect 13737 5661 13771 5695
rect 3893 5593 3927 5627
rect 4353 5593 4387 5627
rect 6009 5593 6043 5627
rect 13829 5593 13863 5627
rect 17141 5593 17175 5627
rect 1409 5525 1443 5559
rect 1685 5525 1719 5559
rect 1961 5525 1995 5559
rect 5825 5525 5859 5559
rect 6837 5525 6871 5559
rect 8401 5525 8435 5559
rect 10977 5525 11011 5559
rect 12081 5525 12115 5559
rect 12633 5525 12667 5559
rect 14105 5525 14139 5559
rect 16405 5525 16439 5559
rect 3249 5321 3283 5355
rect 3525 5321 3559 5355
rect 9505 5321 9539 5355
rect 13277 5321 13311 5355
rect 15025 5321 15059 5355
rect 17049 5321 17083 5355
rect 17969 5321 18003 5355
rect 18797 5321 18831 5355
rect 1777 5253 1811 5287
rect 5181 5253 5215 5287
rect 5457 5253 5491 5287
rect 6009 5253 6043 5287
rect 8033 5253 8067 5287
rect 11805 5253 11839 5287
rect 1501 5185 1535 5219
rect 3617 5185 3651 5219
rect 3801 5185 3835 5219
rect 4813 5185 4847 5219
rect 4967 5185 5001 5219
rect 7021 5185 7055 5219
rect 7297 5185 7331 5219
rect 7451 5185 7485 5219
rect 14657 5185 14691 5219
rect 14750 5185 14784 5219
rect 15393 5185 15427 5219
rect 17325 5185 17359 5219
rect 17417 5185 17451 5219
rect 17509 5185 17543 5219
rect 17693 5185 17727 5219
rect 17877 5185 17911 5219
rect 18613 5185 18647 5219
rect 5365 5117 5399 5151
rect 7757 5117 7791 5151
rect 11069 5117 11103 5151
rect 11345 5117 11379 5151
rect 11529 5117 11563 5151
rect 3341 5049 3375 5083
rect 7113 4981 7147 5015
rect 7481 4981 7515 5015
rect 9597 4981 9631 5015
rect 15485 4981 15519 5015
rect 2605 4777 2639 4811
rect 3939 4777 3973 4811
rect 7757 4777 7791 4811
rect 9597 4777 9631 4811
rect 11161 4777 11195 4811
rect 16405 4777 16439 4811
rect 2881 4641 2915 4675
rect 4077 4641 4111 4675
rect 11989 4641 12023 4675
rect 12173 4641 12207 4675
rect 16129 4641 16163 4675
rect 1409 4573 1443 4607
rect 2513 4573 2547 4607
rect 2789 4573 2823 4607
rect 3801 4573 3835 4607
rect 4261 4573 4295 4607
rect 6009 4573 6043 4607
rect 9689 4573 9723 4607
rect 10701 4573 10735 4607
rect 10977 4573 11011 4607
rect 11253 4573 11287 4607
rect 11437 4573 11471 4607
rect 14381 4573 14415 4607
rect 16221 4573 16255 4607
rect 16314 4573 16348 4607
rect 18091 4573 18125 4607
rect 18245 4573 18279 4607
rect 18613 4573 18647 4607
rect 2237 4505 2271 4539
rect 6285 4505 6319 4539
rect 14657 4505 14691 4539
rect 4169 4437 4203 4471
rect 10793 4437 10827 4471
rect 11253 4437 11287 4471
rect 12633 4437 12667 4471
rect 17877 4437 17911 4471
rect 18797 4437 18831 4471
rect 5273 4233 5307 4267
rect 1685 4097 1719 4131
rect 2053 4097 2087 4131
rect 3249 4097 3283 4131
rect 3433 4097 3467 4131
rect 5457 4097 5491 4131
rect 5549 4097 5583 4131
rect 6653 4097 6687 4131
rect 6837 4097 6871 4131
rect 6929 4097 6963 4131
rect 7205 4097 7239 4131
rect 7757 4097 7791 4131
rect 8891 4097 8925 4131
rect 9045 4097 9079 4131
rect 12541 4097 12575 4131
rect 12633 4097 12667 4131
rect 12725 4097 12759 4131
rect 12909 4097 12943 4131
rect 13461 4097 13495 4131
rect 15209 4097 15243 4131
rect 15393 4097 15427 4131
rect 15485 4097 15519 4131
rect 16037 4097 16071 4131
rect 1593 4029 1627 4063
rect 3525 4029 3559 4063
rect 3801 4029 3835 4063
rect 7573 4029 7607 4063
rect 15853 4029 15887 4063
rect 17049 4029 17083 4063
rect 17325 4029 17359 4063
rect 2237 3961 2271 3995
rect 3341 3961 3375 3995
rect 8677 3961 8711 3995
rect 2053 3893 2087 3927
rect 6469 3893 6503 3927
rect 7113 3893 7147 3927
rect 8217 3893 8251 3927
rect 12265 3893 12299 3927
rect 13369 3893 13403 3927
rect 15025 3893 15059 3927
rect 16497 3893 16531 3927
rect 18797 3893 18831 3927
rect 2697 3689 2731 3723
rect 7481 3689 7515 3723
rect 10701 3689 10735 3723
rect 11897 3689 11931 3723
rect 12430 3689 12464 3723
rect 15853 3689 15887 3723
rect 16037 3689 16071 3723
rect 17233 3689 17267 3723
rect 18337 3689 18371 3723
rect 18521 3689 18555 3723
rect 5549 3553 5583 3587
rect 5825 3553 5859 3587
rect 7297 3553 7331 3587
rect 8953 3553 8987 3587
rect 12173 3553 12207 3587
rect 14105 3553 14139 3587
rect 1409 3485 1443 3519
rect 3801 3485 3835 3519
rect 7389 3485 7423 3519
rect 7573 3485 7607 3519
rect 8125 3485 8159 3519
rect 8309 3485 8343 3519
rect 8401 3485 8435 3519
rect 8493 3485 8527 3519
rect 11927 3485 11961 3519
rect 12081 3485 12115 3519
rect 15945 3485 15979 3519
rect 16129 3485 16163 3519
rect 17509 3485 17543 3519
rect 17601 3485 17635 3519
rect 17693 3485 17727 3519
rect 17877 3485 17911 3519
rect 18153 3485 18187 3519
rect 18429 3485 18463 3519
rect 8769 3417 8803 3451
rect 9229 3417 9263 3451
rect 14381 3417 14415 3451
rect 3893 3349 3927 3383
rect 13921 3349 13955 3383
rect 1593 3145 1627 3179
rect 9781 3145 9815 3179
rect 15669 3145 15703 3179
rect 15853 3145 15887 3179
rect 3985 3077 4019 3111
rect 5641 3077 5675 3111
rect 6837 3077 6871 3111
rect 10885 3077 10919 3111
rect 15485 3077 15519 3111
rect 1409 3009 1443 3043
rect 3709 3009 3743 3043
rect 5733 3009 5767 3043
rect 5825 3009 5859 3043
rect 6469 3009 6503 3043
rect 7113 3009 7147 3043
rect 8953 3009 8987 3043
rect 9689 3009 9723 3043
rect 10057 3009 10091 3043
rect 11153 3009 11187 3043
rect 11529 3009 11563 3043
rect 13369 3009 13403 3043
rect 13737 3009 13771 3043
rect 15945 3009 15979 3043
rect 16670 3009 16704 3043
rect 18521 3009 18555 3043
rect 5457 2941 5491 2975
rect 7389 2941 7423 2975
rect 8861 2941 8895 2975
rect 10517 2941 10551 2975
rect 11805 2941 11839 2975
rect 13277 2941 13311 2975
rect 15117 2941 15151 2975
rect 16957 2941 16991 2975
rect 18429 2941 18463 2975
rect 7021 2873 7055 2907
rect 11069 2873 11103 2907
rect 6009 2805 6043 2839
rect 6837 2805 6871 2839
rect 9137 2805 9171 2839
rect 10241 2805 10275 2839
rect 10885 2805 10919 2839
rect 11345 2805 11379 2839
rect 13553 2805 13587 2839
rect 13921 2805 13955 2839
rect 15485 2805 15519 2839
rect 18705 2805 18739 2839
rect 6101 2601 6135 2635
rect 7205 2601 7239 2635
rect 8217 2601 8251 2635
rect 11069 2601 11103 2635
rect 11805 2601 11839 2635
rect 15577 2601 15611 2635
rect 17325 2601 17359 2635
rect 17509 2601 17543 2635
rect 17785 2601 17819 2635
rect 18061 2601 18095 2635
rect 18797 2601 18831 2635
rect 8033 2533 8067 2567
rect 11989 2533 12023 2567
rect 18337 2533 18371 2567
rect 5917 2397 5951 2431
rect 6745 2397 6779 2431
rect 7389 2397 7423 2431
rect 7849 2397 7883 2431
rect 8125 2397 8159 2431
rect 9321 2397 9355 2431
rect 10609 2397 10643 2431
rect 11253 2397 11287 2431
rect 11713 2397 11747 2431
rect 12173 2397 12207 2431
rect 12357 2397 12391 2431
rect 13829 2397 13863 2431
rect 14473 2397 14507 2431
rect 15761 2397 15795 2431
rect 17233 2397 17267 2431
rect 17693 2397 17727 2431
rect 17969 2397 18003 2431
rect 18245 2397 18279 2431
rect 18521 2397 18555 2431
rect 18613 2397 18647 2431
rect 6561 2261 6595 2295
rect 9137 2261 9171 2295
rect 10425 2261 10459 2295
rect 12541 2261 12575 2295
rect 13645 2261 13679 2295
rect 14289 2261 14323 2295
<< metal1 >>
rect 1104 20154 19136 20176
rect 1104 20102 2350 20154
rect 2402 20102 2414 20154
rect 2466 20102 2478 20154
rect 2530 20102 2542 20154
rect 2594 20102 2606 20154
rect 2658 20102 19136 20154
rect 1104 20080 19136 20102
rect 5258 20000 5264 20052
rect 5316 20000 5322 20052
rect 8478 20000 8484 20052
rect 8536 20000 8542 20052
rect 9766 20000 9772 20052
rect 9824 20000 9830 20052
rect 10870 20000 10876 20052
rect 10928 20040 10934 20052
rect 11057 20043 11115 20049
rect 11057 20040 11069 20043
rect 10928 20012 11069 20040
rect 10928 20000 10934 20012
rect 11057 20009 11069 20012
rect 11103 20009 11115 20043
rect 11057 20003 11115 20009
rect 11698 20000 11704 20052
rect 11756 20000 11762 20052
rect 12986 20000 12992 20052
rect 13044 20000 13050 20052
rect 14274 20000 14280 20052
rect 14332 20000 14338 20052
rect 17494 20000 17500 20052
rect 17552 20000 17558 20052
rect 17770 20000 17776 20052
rect 17828 20000 17834 20052
rect 10597 19975 10655 19981
rect 10597 19941 10609 19975
rect 10643 19941 10655 19975
rect 10597 19935 10655 19941
rect 18417 19975 18475 19981
rect 18417 19941 18429 19975
rect 18463 19941 18475 19975
rect 18417 19935 18475 19941
rect 10612 19904 10640 19935
rect 18432 19904 18460 19935
rect 10612 19876 11284 19904
rect 4890 19796 4896 19848
rect 4948 19836 4954 19848
rect 5445 19839 5503 19845
rect 5445 19836 5457 19839
rect 4948 19808 5457 19836
rect 4948 19796 4954 19808
rect 5445 19805 5457 19808
rect 5491 19805 5503 19839
rect 5445 19799 5503 19805
rect 5902 19796 5908 19848
rect 5960 19796 5966 19848
rect 6730 19796 6736 19848
rect 6788 19796 6794 19848
rect 7190 19796 7196 19848
rect 7248 19796 7254 19848
rect 8662 19796 8668 19848
rect 8720 19796 8726 19848
rect 9155 19839 9213 19845
rect 9155 19836 9167 19839
rect 8772 19808 9167 19836
rect 8772 19768 8800 19808
rect 9155 19805 9167 19808
rect 9201 19805 9213 19839
rect 9155 19799 9213 19805
rect 9309 19839 9367 19845
rect 9309 19805 9321 19839
rect 9355 19805 9367 19839
rect 9309 19799 9367 19805
rect 8404 19740 8800 19768
rect 9324 19768 9352 19799
rect 9950 19796 9956 19848
rect 10008 19796 10014 19848
rect 10413 19839 10471 19845
rect 10413 19805 10425 19839
rect 10459 19805 10471 19839
rect 10413 19799 10471 19805
rect 9490 19768 9496 19780
rect 9324 19740 9496 19768
rect 8404 19712 8432 19740
rect 9490 19728 9496 19740
rect 9548 19768 9554 19780
rect 10428 19768 10456 19799
rect 10594 19796 10600 19848
rect 10652 19836 10658 19848
rect 11256 19845 11284 19876
rect 17328 19876 18460 19904
rect 10873 19839 10931 19845
rect 10873 19836 10885 19839
rect 10652 19808 10885 19836
rect 10652 19796 10658 19808
rect 10873 19805 10885 19808
rect 10919 19805 10931 19839
rect 10873 19799 10931 19805
rect 11241 19839 11299 19845
rect 11241 19805 11253 19839
rect 11287 19805 11299 19839
rect 11241 19799 11299 19805
rect 11698 19796 11704 19848
rect 11756 19836 11762 19848
rect 11885 19839 11943 19845
rect 11885 19836 11897 19839
rect 11756 19808 11897 19836
rect 11756 19796 11762 19808
rect 11885 19805 11897 19808
rect 11931 19805 11943 19839
rect 11885 19799 11943 19805
rect 13173 19839 13231 19845
rect 13173 19805 13185 19839
rect 13219 19836 13231 19839
rect 13262 19836 13268 19848
rect 13219 19808 13268 19836
rect 13219 19805 13231 19808
rect 13173 19799 13231 19805
rect 13262 19796 13268 19808
rect 13320 19796 13326 19848
rect 13722 19796 13728 19848
rect 13780 19836 13786 19848
rect 13817 19839 13875 19845
rect 13817 19836 13829 19839
rect 13780 19808 13829 19836
rect 13780 19796 13786 19808
rect 13817 19805 13829 19808
rect 13863 19805 13875 19839
rect 13817 19799 13875 19805
rect 14458 19796 14464 19848
rect 14516 19796 14522 19848
rect 14918 19796 14924 19848
rect 14976 19796 14982 19848
rect 16206 19796 16212 19848
rect 16264 19796 16270 19848
rect 17328 19845 17356 19876
rect 17313 19839 17371 19845
rect 17313 19805 17325 19839
rect 17359 19805 17371 19839
rect 17313 19799 17371 19805
rect 17589 19839 17647 19845
rect 17589 19805 17601 19839
rect 17635 19805 17647 19839
rect 17589 19799 17647 19805
rect 9548 19740 10456 19768
rect 17604 19768 17632 19799
rect 17862 19796 17868 19848
rect 17920 19796 17926 19848
rect 18230 19796 18236 19848
rect 18288 19836 18294 19848
rect 18325 19839 18383 19845
rect 18325 19836 18337 19839
rect 18288 19808 18337 19836
rect 18288 19796 18294 19808
rect 18325 19805 18337 19808
rect 18371 19805 18383 19839
rect 18325 19799 18383 19805
rect 18506 19796 18512 19848
rect 18564 19836 18570 19848
rect 18601 19839 18659 19845
rect 18601 19836 18613 19839
rect 18564 19808 18613 19836
rect 18564 19796 18570 19808
rect 18601 19805 18613 19808
rect 18647 19805 18659 19839
rect 18601 19799 18659 19805
rect 17604 19740 18184 19768
rect 9548 19728 9554 19740
rect 5718 19660 5724 19712
rect 5776 19700 5782 19712
rect 6089 19703 6147 19709
rect 6089 19700 6101 19703
rect 5776 19672 6101 19700
rect 5776 19660 5782 19672
rect 6089 19669 6101 19672
rect 6135 19669 6147 19703
rect 6089 19663 6147 19669
rect 6546 19660 6552 19712
rect 6604 19660 6610 19712
rect 7377 19703 7435 19709
rect 7377 19669 7389 19703
rect 7423 19700 7435 19703
rect 8386 19700 8392 19712
rect 7423 19672 8392 19700
rect 7423 19669 7435 19672
rect 7377 19663 7435 19669
rect 8386 19660 8392 19672
rect 8444 19660 8450 19712
rect 8941 19703 8999 19709
rect 8941 19669 8953 19703
rect 8987 19700 8999 19703
rect 9398 19700 9404 19712
rect 8987 19672 9404 19700
rect 8987 19669 8999 19672
rect 8941 19663 8999 19669
rect 9398 19660 9404 19672
rect 9456 19660 9462 19712
rect 10502 19660 10508 19712
rect 10560 19700 10566 19712
rect 10689 19703 10747 19709
rect 10689 19700 10701 19703
rect 10560 19672 10701 19700
rect 10560 19660 10566 19672
rect 10689 19669 10701 19672
rect 10735 19669 10747 19703
rect 10689 19663 10747 19669
rect 12894 19660 12900 19712
rect 12952 19700 12958 19712
rect 13633 19703 13691 19709
rect 13633 19700 13645 19703
rect 12952 19672 13645 19700
rect 12952 19660 12958 19672
rect 13633 19669 13645 19672
rect 13679 19669 13691 19703
rect 13633 19663 13691 19669
rect 14918 19660 14924 19712
rect 14976 19700 14982 19712
rect 15105 19703 15163 19709
rect 15105 19700 15117 19703
rect 14976 19672 15117 19700
rect 14976 19660 14982 19672
rect 15105 19669 15117 19672
rect 15151 19669 15163 19703
rect 15105 19663 15163 19669
rect 16390 19660 16396 19712
rect 16448 19660 16454 19712
rect 18046 19660 18052 19712
rect 18104 19660 18110 19712
rect 18156 19709 18184 19740
rect 18141 19703 18199 19709
rect 18141 19669 18153 19703
rect 18187 19669 18199 19703
rect 18141 19663 18199 19669
rect 1104 19610 19136 19632
rect 1104 19558 3010 19610
rect 3062 19558 3074 19610
rect 3126 19558 3138 19610
rect 3190 19558 3202 19610
rect 3254 19558 3266 19610
rect 3318 19558 19136 19610
rect 1104 19536 19136 19558
rect 4433 19499 4491 19505
rect 4433 19465 4445 19499
rect 4479 19465 4491 19499
rect 4433 19459 4491 19465
rect 2866 19428 2872 19440
rect 2700 19400 2872 19428
rect 2700 19369 2728 19400
rect 2866 19388 2872 19400
rect 2924 19388 2930 19440
rect 3970 19388 3976 19440
rect 4028 19388 4034 19440
rect 2685 19363 2743 19369
rect 2685 19329 2697 19363
rect 2731 19329 2743 19363
rect 4448 19360 4476 19459
rect 4890 19456 4896 19508
rect 4948 19456 4954 19508
rect 6546 19456 6552 19508
rect 6604 19456 6610 19508
rect 9490 19456 9496 19508
rect 9548 19456 9554 19508
rect 11333 19499 11391 19505
rect 11333 19465 11345 19499
rect 11379 19465 11391 19499
rect 11333 19459 11391 19465
rect 5644 19400 6040 19428
rect 5644 19369 5672 19400
rect 4709 19363 4767 19369
rect 4709 19360 4721 19363
rect 4448 19332 4721 19360
rect 2685 19323 2743 19329
rect 4709 19329 4721 19332
rect 4755 19329 4767 19363
rect 4709 19323 4767 19329
rect 5629 19363 5687 19369
rect 5629 19329 5641 19363
rect 5675 19329 5687 19363
rect 5629 19323 5687 19329
rect 5718 19320 5724 19372
rect 5776 19320 5782 19372
rect 5902 19320 5908 19372
rect 5960 19320 5966 19372
rect 6012 19360 6040 19400
rect 6638 19388 6644 19440
rect 6696 19428 6702 19440
rect 9306 19428 9312 19440
rect 6696 19400 7788 19428
rect 9246 19400 9312 19428
rect 6696 19388 6702 19400
rect 6730 19360 6736 19372
rect 6012 19332 6736 19360
rect 6730 19320 6736 19332
rect 6788 19360 6794 19372
rect 7760 19369 7788 19400
rect 9306 19388 9312 19400
rect 9364 19388 9370 19440
rect 11348 19428 11376 19459
rect 11698 19456 11704 19508
rect 11756 19456 11762 19508
rect 13262 19456 13268 19508
rect 13320 19456 13326 19508
rect 13817 19499 13875 19505
rect 13817 19465 13829 19499
rect 13863 19496 13875 19499
rect 14458 19496 14464 19508
rect 13863 19468 14464 19496
rect 13863 19465 13875 19468
rect 13817 19459 13875 19465
rect 14458 19456 14464 19468
rect 14516 19456 14522 19508
rect 14918 19456 14924 19508
rect 14976 19456 14982 19508
rect 17862 19456 17868 19508
rect 17920 19496 17926 19508
rect 18509 19499 18567 19505
rect 18509 19496 18521 19499
rect 17920 19468 18521 19496
rect 17920 19456 17926 19468
rect 18509 19465 18521 19468
rect 18555 19465 18567 19499
rect 18509 19459 18567 19465
rect 11348 19400 13124 19428
rect 7193 19363 7251 19369
rect 7193 19360 7205 19363
rect 6788 19332 7205 19360
rect 6788 19320 6794 19332
rect 7193 19329 7205 19332
rect 7239 19329 7251 19363
rect 7193 19323 7251 19329
rect 7745 19363 7803 19369
rect 7745 19329 7757 19363
rect 7791 19329 7803 19363
rect 7745 19323 7803 19329
rect 9582 19320 9588 19372
rect 9640 19320 9646 19372
rect 10962 19320 10968 19372
rect 11020 19320 11026 19372
rect 11514 19320 11520 19372
rect 11572 19320 11578 19372
rect 12894 19360 12900 19372
rect 12855 19332 12900 19360
rect 12894 19320 12900 19332
rect 12952 19320 12958 19372
rect 13096 19369 13124 19400
rect 16942 19388 16948 19440
rect 17000 19428 17006 19440
rect 17000 19400 17434 19428
rect 17000 19388 17006 19400
rect 12989 19363 13047 19369
rect 12989 19329 13001 19363
rect 13035 19329 13047 19363
rect 12989 19323 13047 19329
rect 13081 19363 13139 19369
rect 13081 19329 13093 19363
rect 13127 19329 13139 19363
rect 13081 19323 13139 19329
rect 2961 19295 3019 19301
rect 2961 19292 2973 19295
rect 2700 19264 2973 19292
rect 2700 19236 2728 19264
rect 2961 19261 2973 19264
rect 3007 19261 3019 19295
rect 2961 19255 3019 19261
rect 8021 19295 8079 19301
rect 8021 19261 8033 19295
rect 8067 19292 8079 19295
rect 8754 19292 8760 19304
rect 8067 19264 8760 19292
rect 8067 19261 8079 19264
rect 8021 19255 8079 19261
rect 8754 19252 8760 19264
rect 8812 19252 8818 19304
rect 9861 19295 9919 19301
rect 9861 19261 9873 19295
rect 9907 19292 9919 19295
rect 10594 19292 10600 19304
rect 9907 19264 10600 19292
rect 9907 19261 9919 19264
rect 9861 19255 9919 19261
rect 10594 19252 10600 19264
rect 10652 19252 10658 19304
rect 13004 19292 13032 19323
rect 13630 19320 13636 19372
rect 13688 19320 13694 19372
rect 15194 19320 15200 19372
rect 15252 19320 15258 19372
rect 15381 19363 15439 19369
rect 15381 19329 15393 19363
rect 15427 19360 15439 19363
rect 16390 19360 16396 19372
rect 15427 19332 16396 19360
rect 15427 19329 15439 19332
rect 15381 19323 15439 19329
rect 13648 19292 13676 19320
rect 15396 19292 15424 19323
rect 16390 19320 16396 19332
rect 16448 19320 16454 19372
rect 18690 19320 18696 19372
rect 18748 19320 18754 19372
rect 13004 19264 13676 19292
rect 14752 19264 15424 19292
rect 2682 19184 2688 19236
rect 2740 19184 2746 19236
rect 5718 19184 5724 19236
rect 5776 19224 5782 19236
rect 6917 19227 6975 19233
rect 5776 19196 6592 19224
rect 5776 19184 5782 19196
rect 5537 19159 5595 19165
rect 5537 19125 5549 19159
rect 5583 19156 5595 19159
rect 5626 19156 5632 19168
rect 5583 19128 5632 19156
rect 5583 19125 5595 19128
rect 5537 19119 5595 19125
rect 5626 19116 5632 19128
rect 5684 19116 5690 19168
rect 5810 19116 5816 19168
rect 5868 19116 5874 19168
rect 6365 19159 6423 19165
rect 6365 19125 6377 19159
rect 6411 19156 6423 19159
rect 6454 19156 6460 19168
rect 6411 19128 6460 19156
rect 6411 19125 6423 19128
rect 6365 19119 6423 19125
rect 6454 19116 6460 19128
rect 6512 19116 6518 19168
rect 6564 19165 6592 19196
rect 6917 19193 6929 19227
rect 6963 19224 6975 19227
rect 14553 19227 14611 19233
rect 14553 19224 14565 19227
rect 6963 19196 7420 19224
rect 6963 19193 6975 19196
rect 6917 19187 6975 19193
rect 6549 19159 6607 19165
rect 6549 19125 6561 19159
rect 6595 19156 6607 19159
rect 6822 19156 6828 19168
rect 6595 19128 6828 19156
rect 6595 19125 6607 19128
rect 6549 19119 6607 19125
rect 6822 19116 6828 19128
rect 6880 19116 6886 19168
rect 7190 19116 7196 19168
rect 7248 19156 7254 19168
rect 7285 19159 7343 19165
rect 7285 19156 7297 19159
rect 7248 19128 7297 19156
rect 7248 19116 7254 19128
rect 7285 19125 7297 19128
rect 7331 19125 7343 19159
rect 7392 19156 7420 19196
rect 12406 19196 14565 19224
rect 10226 19156 10232 19168
rect 7392 19128 10232 19156
rect 7285 19119 7343 19125
rect 10226 19116 10232 19128
rect 10284 19156 10290 19168
rect 11790 19156 11796 19168
rect 10284 19128 11796 19156
rect 10284 19116 10290 19128
rect 11790 19116 11796 19128
rect 11848 19156 11854 19168
rect 12406 19156 12434 19196
rect 14553 19193 14565 19196
rect 14599 19193 14611 19227
rect 14553 19187 14611 19193
rect 11848 19128 12434 19156
rect 11848 19116 11854 19128
rect 12710 19116 12716 19168
rect 12768 19156 12774 19168
rect 12805 19159 12863 19165
rect 12805 19156 12817 19159
rect 12768 19128 12817 19156
rect 12768 19116 12774 19128
rect 12805 19125 12817 19128
rect 12851 19125 12863 19159
rect 14752 19156 14780 19264
rect 16666 19252 16672 19304
rect 16724 19252 16730 19304
rect 16945 19295 17003 19301
rect 16945 19292 16957 19295
rect 16776 19264 16957 19292
rect 14826 19184 14832 19236
rect 14884 19224 14890 19236
rect 15105 19227 15163 19233
rect 15105 19224 15117 19227
rect 14884 19196 15117 19224
rect 14884 19184 14890 19196
rect 15105 19193 15117 19196
rect 15151 19224 15163 19227
rect 16776 19224 16804 19264
rect 16945 19261 16957 19264
rect 16991 19261 17003 19295
rect 16945 19255 17003 19261
rect 15151 19196 16804 19224
rect 15151 19193 15163 19196
rect 15105 19187 15163 19193
rect 14921 19159 14979 19165
rect 14921 19156 14933 19159
rect 14752 19128 14933 19156
rect 12805 19119 12863 19125
rect 14921 19125 14933 19128
rect 14967 19125 14979 19159
rect 14921 19119 14979 19125
rect 15286 19116 15292 19168
rect 15344 19116 15350 19168
rect 18414 19116 18420 19168
rect 18472 19116 18478 19168
rect 1104 19066 19136 19088
rect 1104 19014 2350 19066
rect 2402 19014 2414 19066
rect 2466 19014 2478 19066
rect 2530 19014 2542 19066
rect 2594 19014 2606 19066
rect 2658 19014 19136 19066
rect 1104 18992 19136 19014
rect 3881 18955 3939 18961
rect 3881 18921 3893 18955
rect 3927 18952 3939 18955
rect 3970 18952 3976 18964
rect 3927 18924 3976 18952
rect 3927 18921 3939 18924
rect 3881 18915 3939 18921
rect 3970 18912 3976 18924
rect 4028 18912 4034 18964
rect 8205 18955 8263 18961
rect 8205 18921 8217 18955
rect 8251 18952 8263 18955
rect 8662 18952 8668 18964
rect 8251 18924 8668 18952
rect 8251 18921 8263 18924
rect 8205 18915 8263 18921
rect 8662 18912 8668 18924
rect 8720 18912 8726 18964
rect 8754 18912 8760 18964
rect 8812 18952 8818 18964
rect 8941 18955 8999 18961
rect 8941 18952 8953 18955
rect 8812 18924 8953 18952
rect 8812 18912 8818 18924
rect 8941 18921 8953 18924
rect 8987 18921 8999 18955
rect 8941 18915 8999 18921
rect 9306 18912 9312 18964
rect 9364 18952 9370 18964
rect 9769 18955 9827 18961
rect 9769 18952 9781 18955
rect 9364 18924 9781 18952
rect 9364 18912 9370 18924
rect 9769 18921 9781 18924
rect 9815 18921 9827 18955
rect 9769 18915 9827 18921
rect 10505 18955 10563 18961
rect 10505 18921 10517 18955
rect 10551 18921 10563 18955
rect 10505 18915 10563 18921
rect 10137 18887 10195 18893
rect 10137 18853 10149 18887
rect 10183 18884 10195 18887
rect 10226 18884 10232 18896
rect 10183 18856 10232 18884
rect 10183 18853 10195 18856
rect 10137 18847 10195 18853
rect 10226 18844 10232 18856
rect 10284 18844 10290 18896
rect 10520 18884 10548 18915
rect 10594 18912 10600 18964
rect 10652 18952 10658 18964
rect 10689 18955 10747 18961
rect 10689 18952 10701 18955
rect 10652 18924 10701 18952
rect 10652 18912 10658 18924
rect 10689 18921 10701 18924
rect 10735 18921 10747 18955
rect 10689 18915 10747 18921
rect 10962 18912 10968 18964
rect 11020 18952 11026 18964
rect 11609 18955 11667 18961
rect 11609 18952 11621 18955
rect 11020 18924 11621 18952
rect 11020 18912 11026 18924
rect 11609 18921 11621 18924
rect 11655 18921 11667 18955
rect 11609 18915 11667 18921
rect 13630 18912 13636 18964
rect 13688 18952 13694 18964
rect 13725 18955 13783 18961
rect 13725 18952 13737 18955
rect 13688 18924 13737 18952
rect 13688 18912 13694 18924
rect 13725 18921 13737 18924
rect 13771 18921 13783 18955
rect 13725 18915 13783 18921
rect 16942 18912 16948 18964
rect 17000 18912 17006 18964
rect 18046 18912 18052 18964
rect 18104 18912 18110 18964
rect 11698 18884 11704 18896
rect 10520 18856 11704 18884
rect 11698 18844 11704 18856
rect 11756 18844 11762 18896
rect 18141 18887 18199 18893
rect 18141 18853 18153 18887
rect 18187 18853 18199 18887
rect 18141 18847 18199 18853
rect 4341 18819 4399 18825
rect 4341 18816 4353 18819
rect 1780 18788 4353 18816
rect 842 18708 848 18760
rect 900 18748 906 18760
rect 1397 18751 1455 18757
rect 1397 18748 1409 18751
rect 900 18720 1409 18748
rect 900 18708 906 18720
rect 1397 18717 1409 18720
rect 1443 18717 1455 18751
rect 1397 18711 1455 18717
rect 1670 18708 1676 18760
rect 1728 18748 1734 18760
rect 1780 18757 1808 18788
rect 4341 18785 4353 18788
rect 4387 18816 4399 18819
rect 6181 18819 6239 18825
rect 6181 18816 6193 18819
rect 4387 18788 6193 18816
rect 4387 18785 4399 18788
rect 4341 18779 4399 18785
rect 6181 18785 6193 18788
rect 6227 18816 6239 18819
rect 6546 18816 6552 18828
rect 6227 18788 6552 18816
rect 6227 18785 6239 18788
rect 6181 18779 6239 18785
rect 6546 18776 6552 18788
rect 6604 18776 6610 18828
rect 7929 18819 7987 18825
rect 7929 18785 7941 18819
rect 7975 18785 7987 18819
rect 7929 18779 7987 18785
rect 1765 18751 1823 18757
rect 1765 18748 1777 18751
rect 1728 18720 1777 18748
rect 1728 18708 1734 18720
rect 1765 18717 1777 18720
rect 1811 18717 1823 18751
rect 1765 18711 1823 18717
rect 3970 18708 3976 18760
rect 4028 18708 4034 18760
rect 7944 18748 7972 18779
rect 9122 18776 9128 18828
rect 9180 18816 9186 18828
rect 9674 18816 9680 18828
rect 9180 18788 9680 18816
rect 9180 18776 9186 18788
rect 8021 18751 8079 18757
rect 8021 18748 8033 18751
rect 7944 18720 8033 18748
rect 8021 18717 8033 18720
rect 8067 18717 8079 18751
rect 8021 18711 8079 18717
rect 8386 18708 8392 18760
rect 8444 18748 8450 18760
rect 9324 18757 9352 18788
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 11146 18816 11152 18828
rect 9876 18788 11152 18816
rect 9217 18751 9275 18757
rect 9217 18748 9229 18751
rect 8444 18720 9229 18748
rect 8444 18708 8450 18720
rect 9217 18717 9229 18720
rect 9263 18717 9275 18751
rect 9217 18711 9275 18717
rect 9309 18751 9367 18757
rect 9309 18717 9321 18751
rect 9355 18717 9367 18751
rect 9309 18711 9367 18717
rect 9398 18708 9404 18760
rect 9456 18708 9462 18760
rect 9876 18757 9904 18788
rect 11146 18776 11152 18788
rect 11204 18816 11210 18828
rect 11977 18819 12035 18825
rect 11204 18788 11744 18816
rect 11204 18776 11210 18788
rect 11716 18757 11744 18788
rect 11977 18785 11989 18819
rect 12023 18816 12035 18819
rect 12618 18816 12624 18828
rect 12023 18788 12624 18816
rect 12023 18785 12035 18788
rect 11977 18779 12035 18785
rect 12618 18776 12624 18788
rect 12676 18816 12682 18828
rect 14093 18819 14151 18825
rect 14093 18816 14105 18819
rect 12676 18788 14105 18816
rect 12676 18776 12682 18788
rect 14093 18785 14105 18788
rect 14139 18785 14151 18819
rect 14093 18779 14151 18785
rect 9585 18751 9643 18757
rect 9585 18717 9597 18751
rect 9631 18717 9643 18751
rect 9585 18711 9643 18717
rect 9861 18751 9919 18757
rect 9861 18717 9873 18751
rect 9907 18717 9919 18751
rect 9861 18711 9919 18717
rect 11701 18751 11759 18757
rect 11701 18717 11713 18751
rect 11747 18717 11759 18751
rect 11701 18711 11759 18717
rect 2041 18683 2099 18689
rect 2041 18649 2053 18683
rect 2087 18680 2099 18683
rect 2314 18680 2320 18692
rect 2087 18652 2320 18680
rect 2087 18649 2099 18652
rect 2041 18643 2099 18649
rect 2314 18640 2320 18652
rect 2372 18640 2378 18692
rect 3418 18680 3424 18692
rect 3266 18652 3424 18680
rect 3418 18640 3424 18652
rect 3476 18640 3482 18692
rect 4614 18640 4620 18692
rect 4672 18640 4678 18692
rect 5626 18640 5632 18692
rect 5684 18640 5690 18692
rect 6454 18640 6460 18692
rect 6512 18640 6518 18692
rect 7190 18640 7196 18692
rect 7248 18640 7254 18692
rect 1581 18615 1639 18621
rect 1581 18581 1593 18615
rect 1627 18612 1639 18615
rect 1762 18612 1768 18624
rect 1627 18584 1768 18612
rect 1627 18581 1639 18584
rect 1581 18575 1639 18581
rect 1762 18572 1768 18584
rect 1820 18572 1826 18624
rect 3510 18572 3516 18624
rect 3568 18572 3574 18624
rect 5994 18572 6000 18624
rect 6052 18612 6058 18624
rect 6089 18615 6147 18621
rect 6089 18612 6101 18615
rect 6052 18584 6101 18612
rect 6052 18572 6058 18584
rect 6089 18581 6101 18584
rect 6135 18581 6147 18615
rect 6089 18575 6147 18581
rect 7374 18572 7380 18624
rect 7432 18612 7438 18624
rect 9600 18612 9628 18711
rect 16390 18708 16396 18760
rect 16448 18748 16454 18760
rect 16607 18751 16665 18757
rect 16607 18748 16619 18751
rect 16448 18720 16619 18748
rect 16448 18708 16454 18720
rect 16607 18717 16619 18720
rect 16653 18717 16665 18751
rect 16607 18711 16665 18717
rect 16761 18751 16819 18757
rect 16761 18717 16773 18751
rect 16807 18717 16819 18751
rect 16761 18711 16819 18717
rect 10502 18640 10508 18692
rect 10560 18640 10566 18692
rect 12158 18640 12164 18692
rect 12216 18680 12222 18692
rect 12253 18683 12311 18689
rect 12253 18680 12265 18683
rect 12216 18652 12265 18680
rect 12216 18640 12222 18652
rect 12253 18649 12265 18652
rect 12299 18649 12311 18683
rect 12253 18643 12311 18649
rect 12986 18640 12992 18692
rect 13044 18640 13050 18692
rect 14369 18683 14427 18689
rect 14369 18649 14381 18683
rect 14415 18680 14427 18683
rect 14642 18680 14648 18692
rect 14415 18652 14648 18680
rect 14415 18649 14427 18652
rect 14369 18643 14427 18649
rect 14642 18640 14648 18652
rect 14700 18640 14706 18692
rect 15378 18640 15384 18692
rect 15436 18640 15442 18692
rect 16776 18680 16804 18711
rect 16850 18708 16856 18760
rect 16908 18708 16914 18760
rect 17865 18751 17923 18757
rect 17865 18717 17877 18751
rect 17911 18748 17923 18751
rect 18156 18748 18184 18847
rect 18322 18748 18328 18760
rect 17911 18720 18184 18748
rect 18248 18720 18328 18748
rect 17911 18717 17923 18720
rect 17865 18711 17923 18717
rect 18248 18680 18276 18720
rect 18322 18708 18328 18720
rect 18380 18708 18386 18760
rect 18414 18708 18420 18760
rect 18472 18708 18478 18760
rect 16776 18652 18276 18680
rect 11422 18612 11428 18624
rect 7432 18584 11428 18612
rect 7432 18572 7438 18584
rect 11422 18572 11428 18584
rect 11480 18572 11486 18624
rect 15654 18572 15660 18624
rect 15712 18612 15718 18624
rect 15841 18615 15899 18621
rect 15841 18612 15853 18615
rect 15712 18584 15853 18612
rect 15712 18572 15718 18584
rect 15841 18581 15853 18584
rect 15887 18581 15899 18615
rect 15841 18575 15899 18581
rect 16393 18615 16451 18621
rect 16393 18581 16405 18615
rect 16439 18612 16451 18615
rect 16482 18612 16488 18624
rect 16439 18584 16488 18612
rect 16439 18581 16451 18584
rect 16393 18575 16451 18581
rect 16482 18572 16488 18584
rect 16540 18572 16546 18624
rect 18598 18572 18604 18624
rect 18656 18572 18662 18624
rect 1104 18522 19136 18544
rect 1104 18470 3010 18522
rect 3062 18470 3074 18522
rect 3126 18470 3138 18522
rect 3190 18470 3202 18522
rect 3254 18470 3266 18522
rect 3318 18470 19136 18522
rect 1104 18448 19136 18470
rect 1581 18411 1639 18417
rect 1581 18377 1593 18411
rect 1627 18377 1639 18411
rect 1581 18371 1639 18377
rect 1596 18340 1624 18371
rect 1762 18368 1768 18420
rect 1820 18368 1826 18420
rect 2314 18368 2320 18420
rect 2372 18368 2378 18420
rect 2685 18411 2743 18417
rect 2685 18377 2697 18411
rect 2731 18408 2743 18411
rect 2869 18411 2927 18417
rect 2869 18408 2881 18411
rect 2731 18380 2881 18408
rect 2731 18377 2743 18380
rect 2685 18371 2743 18377
rect 2869 18377 2881 18380
rect 2915 18377 2927 18411
rect 2869 18371 2927 18377
rect 3237 18411 3295 18417
rect 3237 18377 3249 18411
rect 3283 18408 3295 18411
rect 3418 18408 3424 18420
rect 3283 18380 3424 18408
rect 3283 18377 3295 18380
rect 3237 18371 3295 18377
rect 3418 18368 3424 18380
rect 3476 18368 3482 18420
rect 4614 18368 4620 18420
rect 4672 18408 4678 18420
rect 5537 18411 5595 18417
rect 5537 18408 5549 18411
rect 4672 18380 5549 18408
rect 4672 18368 4678 18380
rect 5537 18377 5549 18380
rect 5583 18377 5595 18411
rect 5537 18371 5595 18377
rect 5810 18368 5816 18420
rect 5868 18408 5874 18420
rect 5905 18411 5963 18417
rect 5905 18408 5917 18411
rect 5868 18380 5917 18408
rect 5868 18368 5874 18380
rect 5905 18377 5917 18380
rect 5951 18377 5963 18411
rect 5905 18371 5963 18377
rect 6822 18368 6828 18420
rect 6880 18408 6886 18420
rect 9401 18411 9459 18417
rect 6880 18380 7696 18408
rect 6880 18368 6886 18380
rect 1596 18312 2544 18340
rect 2516 18281 2544 18312
rect 2590 18300 2596 18352
rect 2648 18340 2654 18352
rect 6454 18340 6460 18352
rect 2648 18312 3096 18340
rect 2648 18300 2654 18312
rect 2501 18275 2559 18281
rect 2501 18241 2513 18275
rect 2547 18272 2559 18275
rect 2682 18272 2688 18284
rect 2547 18244 2688 18272
rect 2547 18241 2559 18244
rect 2501 18235 2559 18241
rect 2682 18232 2688 18244
rect 2740 18232 2746 18284
rect 2777 18275 2835 18281
rect 2777 18241 2789 18275
rect 2823 18241 2835 18275
rect 2777 18235 2835 18241
rect 2869 18275 2927 18281
rect 2869 18241 2881 18275
rect 2915 18272 2927 18275
rect 2958 18272 2964 18284
rect 2915 18244 2964 18272
rect 2915 18241 2927 18244
rect 2869 18235 2927 18241
rect 2792 18204 2820 18235
rect 2958 18232 2964 18244
rect 3016 18232 3022 18284
rect 3068 18281 3096 18312
rect 5736 18312 6460 18340
rect 3053 18275 3111 18281
rect 3053 18241 3065 18275
rect 3099 18241 3111 18275
rect 3053 18235 3111 18241
rect 3326 18232 3332 18284
rect 3384 18272 3390 18284
rect 3970 18272 3976 18284
rect 3384 18244 3976 18272
rect 3384 18232 3390 18244
rect 3970 18232 3976 18244
rect 4028 18232 4034 18284
rect 5736 18281 5764 18312
rect 6454 18300 6460 18312
rect 6512 18300 6518 18352
rect 7193 18343 7251 18349
rect 7193 18309 7205 18343
rect 7239 18340 7251 18343
rect 7239 18312 7604 18340
rect 7239 18309 7251 18312
rect 7193 18303 7251 18309
rect 7576 18284 7604 18312
rect 5721 18275 5779 18281
rect 5721 18241 5733 18275
rect 5767 18241 5779 18275
rect 5721 18235 5779 18241
rect 5994 18232 6000 18284
rect 6052 18272 6058 18284
rect 6549 18275 6607 18281
rect 6549 18272 6561 18275
rect 6052 18244 6561 18272
rect 6052 18232 6058 18244
rect 6549 18241 6561 18244
rect 6595 18241 6607 18275
rect 7285 18275 7343 18281
rect 7285 18272 7297 18275
rect 6549 18235 6607 18241
rect 6656 18244 7297 18272
rect 3510 18204 3516 18216
rect 2792 18176 3516 18204
rect 3510 18164 3516 18176
rect 3568 18164 3574 18216
rect 5902 18164 5908 18216
rect 5960 18204 5966 18216
rect 6656 18204 6684 18244
rect 7285 18241 7297 18244
rect 7331 18272 7343 18275
rect 7374 18272 7380 18284
rect 7331 18244 7380 18272
rect 7331 18241 7343 18244
rect 7285 18235 7343 18241
rect 7374 18232 7380 18244
rect 7432 18232 7438 18284
rect 7469 18275 7527 18281
rect 7469 18241 7481 18275
rect 7515 18241 7527 18275
rect 7469 18235 7527 18241
rect 5960 18176 6684 18204
rect 5960 18164 5966 18176
rect 6730 18164 6736 18216
rect 6788 18164 6794 18216
rect 7484 18204 7512 18235
rect 7558 18232 7564 18284
rect 7616 18232 7622 18284
rect 7668 18281 7696 18380
rect 9401 18377 9413 18411
rect 9447 18408 9459 18411
rect 9950 18408 9956 18420
rect 9447 18380 9956 18408
rect 9447 18377 9459 18380
rect 9401 18371 9459 18377
rect 9950 18368 9956 18380
rect 10008 18368 10014 18420
rect 12158 18368 12164 18420
rect 12216 18368 12222 18420
rect 12268 18380 12848 18408
rect 11422 18300 11428 18352
rect 11480 18340 11486 18352
rect 12268 18340 12296 18380
rect 11480 18312 12296 18340
rect 11480 18300 11486 18312
rect 7653 18275 7711 18281
rect 7653 18241 7665 18275
rect 7699 18272 7711 18275
rect 8235 18275 8293 18281
rect 8235 18272 8247 18275
rect 7699 18244 8247 18272
rect 7699 18241 7711 18244
rect 7653 18235 7711 18241
rect 8235 18241 8247 18244
rect 8281 18241 8293 18275
rect 8235 18235 8293 18241
rect 8389 18275 8447 18281
rect 8389 18241 8401 18275
rect 8435 18272 8447 18275
rect 9214 18272 9220 18284
rect 8435 18244 9220 18272
rect 8435 18241 8447 18244
rect 8389 18235 8447 18241
rect 9214 18232 9220 18244
rect 9272 18232 9278 18284
rect 12391 18275 12449 18281
rect 12391 18241 12403 18275
rect 12437 18241 12449 18275
rect 12526 18256 12532 18308
rect 12584 18256 12590 18308
rect 12621 18278 12679 18284
rect 12526 18247 12538 18256
rect 12572 18247 12584 18256
rect 12526 18241 12584 18247
rect 12621 18244 12633 18278
rect 12667 18275 12679 18278
rect 12710 18275 12716 18284
rect 12667 18247 12716 18275
rect 12667 18244 12679 18247
rect 12391 18235 12449 18241
rect 12621 18238 12679 18244
rect 8021 18207 8079 18213
rect 8021 18204 8033 18207
rect 7484 18176 8033 18204
rect 8021 18173 8033 18176
rect 8067 18173 8079 18207
rect 8021 18167 8079 18173
rect 11698 18164 11704 18216
rect 11756 18204 11762 18216
rect 12406 18204 12434 18235
rect 12710 18232 12716 18247
rect 12768 18232 12774 18284
rect 12820 18281 12848 18380
rect 12986 18368 12992 18420
rect 13044 18408 13050 18420
rect 13081 18411 13139 18417
rect 13081 18408 13093 18411
rect 13044 18380 13093 18408
rect 13044 18368 13050 18380
rect 13081 18377 13093 18380
rect 13127 18377 13139 18411
rect 13081 18371 13139 18377
rect 14642 18368 14648 18420
rect 14700 18368 14706 18420
rect 15013 18411 15071 18417
rect 15013 18377 15025 18411
rect 15059 18408 15071 18411
rect 15286 18408 15292 18420
rect 15059 18380 15292 18408
rect 15059 18377 15071 18380
rect 15013 18371 15071 18377
rect 15286 18368 15292 18380
rect 15344 18368 15350 18420
rect 18322 18368 18328 18420
rect 18380 18408 18386 18420
rect 18417 18411 18475 18417
rect 18417 18408 18429 18411
rect 18380 18380 18429 18408
rect 18380 18368 18386 18380
rect 18417 18377 18429 18380
rect 18463 18377 18475 18411
rect 18417 18371 18475 18377
rect 18782 18368 18788 18420
rect 18840 18368 18846 18420
rect 13004 18312 15424 18340
rect 13004 18281 13032 18312
rect 12805 18275 12863 18281
rect 12805 18241 12817 18275
rect 12851 18241 12863 18275
rect 12805 18235 12863 18241
rect 12989 18275 13047 18281
rect 12989 18241 13001 18275
rect 13035 18241 13047 18275
rect 12989 18235 13047 18241
rect 12894 18204 12900 18216
rect 11756 18176 12900 18204
rect 11756 18164 11762 18176
rect 12894 18164 12900 18176
rect 12952 18164 12958 18216
rect 1946 18096 1952 18148
rect 2004 18136 2010 18148
rect 2133 18139 2191 18145
rect 2133 18136 2145 18139
rect 2004 18108 2145 18136
rect 2004 18096 2010 18108
rect 2133 18105 2145 18108
rect 2179 18105 2191 18139
rect 2133 18099 2191 18105
rect 2774 18096 2780 18148
rect 2832 18136 2838 18148
rect 3326 18136 3332 18148
rect 2832 18108 3332 18136
rect 2832 18096 2838 18108
rect 3326 18096 3332 18108
rect 3384 18096 3390 18148
rect 11146 18096 11152 18148
rect 11204 18136 11210 18148
rect 12710 18136 12716 18148
rect 11204 18108 12716 18136
rect 11204 18096 11210 18108
rect 12710 18096 12716 18108
rect 12768 18136 12774 18148
rect 13004 18136 13032 18235
rect 14826 18232 14832 18284
rect 14884 18232 14890 18284
rect 15396 18281 15424 18312
rect 17678 18300 17684 18352
rect 17736 18300 17742 18352
rect 15105 18275 15163 18281
rect 15105 18241 15117 18275
rect 15151 18241 15163 18275
rect 15105 18235 15163 18241
rect 15381 18275 15439 18281
rect 15381 18241 15393 18275
rect 15427 18241 15439 18275
rect 15381 18235 15439 18241
rect 15565 18275 15623 18281
rect 15565 18241 15577 18275
rect 15611 18272 15623 18275
rect 15654 18272 15660 18284
rect 15611 18244 15660 18272
rect 15611 18241 15623 18244
rect 15565 18235 15623 18241
rect 15120 18204 15148 18235
rect 15580 18204 15608 18235
rect 15654 18232 15660 18244
rect 15712 18232 15718 18284
rect 18598 18232 18604 18284
rect 18656 18232 18662 18284
rect 15120 18176 15608 18204
rect 15746 18164 15752 18216
rect 15804 18164 15810 18216
rect 15838 18164 15844 18216
rect 15896 18204 15902 18216
rect 16666 18204 16672 18216
rect 15896 18176 16672 18204
rect 15896 18164 15902 18176
rect 16666 18164 16672 18176
rect 16724 18164 16730 18216
rect 16942 18164 16948 18216
rect 17000 18164 17006 18216
rect 12768 18108 13032 18136
rect 15289 18139 15347 18145
rect 12768 18096 12774 18108
rect 15289 18105 15301 18139
rect 15335 18136 15347 18139
rect 15378 18136 15384 18148
rect 15335 18108 15384 18136
rect 15335 18105 15347 18108
rect 15289 18099 15347 18105
rect 15378 18096 15384 18108
rect 15436 18096 15442 18148
rect 1578 18028 1584 18080
rect 1636 18068 1642 18080
rect 1765 18071 1823 18077
rect 1765 18068 1777 18071
rect 1636 18040 1777 18068
rect 1636 18028 1642 18040
rect 1765 18037 1777 18040
rect 1811 18068 1823 18071
rect 2222 18068 2228 18080
rect 1811 18040 2228 18068
rect 1811 18037 1823 18040
rect 1765 18031 1823 18037
rect 2222 18028 2228 18040
rect 2280 18068 2286 18080
rect 2590 18068 2596 18080
rect 2280 18040 2596 18068
rect 2280 18028 2286 18040
rect 2590 18028 2596 18040
rect 2648 18028 2654 18080
rect 2958 18028 2964 18080
rect 3016 18068 3022 18080
rect 3418 18068 3424 18080
rect 3016 18040 3424 18068
rect 3016 18028 3022 18040
rect 3418 18028 3424 18040
rect 3476 18068 3482 18080
rect 5902 18068 5908 18080
rect 3476 18040 5908 18068
rect 3476 18028 3482 18040
rect 5902 18028 5908 18040
rect 5960 18028 5966 18080
rect 7926 18028 7932 18080
rect 7984 18028 7990 18080
rect 16209 18071 16267 18077
rect 16209 18037 16221 18071
rect 16255 18068 16267 18071
rect 16574 18068 16580 18080
rect 16255 18040 16580 18068
rect 16255 18037 16267 18040
rect 16209 18031 16267 18037
rect 16574 18028 16580 18040
rect 16632 18028 16638 18080
rect 1104 17978 19136 18000
rect 1104 17926 2350 17978
rect 2402 17926 2414 17978
rect 2466 17926 2478 17978
rect 2530 17926 2542 17978
rect 2594 17926 2606 17978
rect 2658 17926 19136 17978
rect 1104 17904 19136 17926
rect 1578 17824 1584 17876
rect 1636 17824 1642 17876
rect 12342 17824 12348 17876
rect 12400 17824 12406 17876
rect 16942 17824 16948 17876
rect 17000 17824 17006 17876
rect 17678 17824 17684 17876
rect 17736 17824 17742 17876
rect 6730 17756 6736 17808
rect 6788 17756 6794 17808
rect 11330 17728 11336 17740
rect 10888 17700 11336 17728
rect 842 17620 848 17672
rect 900 17660 906 17672
rect 1397 17663 1455 17669
rect 1397 17660 1409 17663
rect 900 17632 1409 17660
rect 900 17620 906 17632
rect 1397 17629 1409 17632
rect 1443 17629 1455 17663
rect 1397 17623 1455 17629
rect 6362 17620 6368 17672
rect 6420 17620 6426 17672
rect 6454 17620 6460 17672
rect 6512 17620 6518 17672
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17660 8631 17663
rect 8662 17660 8668 17672
rect 8619 17632 8668 17660
rect 8619 17629 8631 17632
rect 8573 17623 8631 17629
rect 8662 17620 8668 17632
rect 8720 17620 8726 17672
rect 10594 17620 10600 17672
rect 10652 17620 10658 17672
rect 10888 17669 10916 17700
rect 11330 17688 11336 17700
rect 11388 17728 11394 17740
rect 11793 17731 11851 17737
rect 11793 17728 11805 17731
rect 11388 17700 11805 17728
rect 11388 17688 11394 17700
rect 11793 17697 11805 17700
rect 11839 17697 11851 17731
rect 11793 17691 11851 17697
rect 15565 17731 15623 17737
rect 15565 17697 15577 17731
rect 15611 17728 15623 17731
rect 16390 17728 16396 17740
rect 15611 17700 16396 17728
rect 15611 17697 15623 17700
rect 15565 17691 15623 17697
rect 16390 17688 16396 17700
rect 16448 17728 16454 17740
rect 16448 17700 16712 17728
rect 16448 17688 16454 17700
rect 10873 17663 10931 17669
rect 10873 17629 10885 17663
rect 10919 17629 10931 17663
rect 10873 17623 10931 17629
rect 11146 17620 11152 17672
rect 11204 17620 11210 17672
rect 11882 17620 11888 17672
rect 11940 17660 11946 17672
rect 11977 17663 12035 17669
rect 11977 17660 11989 17663
rect 11940 17632 11989 17660
rect 11940 17620 11946 17632
rect 11977 17629 11989 17632
rect 12023 17629 12035 17663
rect 11977 17623 12035 17629
rect 15838 17620 15844 17672
rect 15896 17620 15902 17672
rect 16301 17663 16359 17669
rect 16301 17629 16313 17663
rect 16347 17629 16359 17663
rect 16301 17623 16359 17629
rect 14826 17552 14832 17604
rect 14884 17552 14890 17604
rect 15286 17552 15292 17604
rect 15344 17592 15350 17604
rect 16316 17592 16344 17623
rect 16482 17620 16488 17672
rect 16540 17620 16546 17672
rect 16574 17620 16580 17672
rect 16632 17620 16638 17672
rect 16684 17669 16712 17700
rect 16669 17663 16727 17669
rect 16669 17629 16681 17663
rect 16715 17629 16727 17663
rect 16669 17623 16727 17629
rect 16850 17620 16856 17672
rect 16908 17660 16914 17672
rect 17589 17663 17647 17669
rect 17589 17660 17601 17663
rect 16908 17632 17601 17660
rect 16908 17620 16914 17632
rect 17589 17629 17601 17632
rect 17635 17660 17647 17663
rect 17862 17660 17868 17672
rect 17635 17632 17868 17660
rect 17635 17629 17647 17632
rect 17589 17623 17647 17629
rect 17862 17620 17868 17632
rect 17920 17620 17926 17672
rect 18782 17620 18788 17672
rect 18840 17620 18846 17672
rect 17770 17592 17776 17604
rect 15344 17564 17776 17592
rect 15344 17552 15350 17564
rect 17770 17552 17776 17564
rect 17828 17552 17834 17604
rect 8570 17484 8576 17536
rect 8628 17524 8634 17536
rect 8665 17527 8723 17533
rect 8665 17524 8677 17527
rect 8628 17496 8677 17524
rect 8628 17484 8634 17496
rect 8665 17493 8677 17496
rect 8711 17493 8723 17527
rect 8665 17487 8723 17493
rect 9858 17484 9864 17536
rect 9916 17524 9922 17536
rect 10413 17527 10471 17533
rect 10413 17524 10425 17527
rect 9916 17496 10425 17524
rect 9916 17484 9922 17496
rect 10413 17493 10425 17496
rect 10459 17493 10471 17527
rect 10413 17487 10471 17493
rect 10778 17484 10784 17536
rect 10836 17484 10842 17536
rect 10870 17484 10876 17536
rect 10928 17524 10934 17536
rect 11057 17527 11115 17533
rect 11057 17524 11069 17527
rect 10928 17496 11069 17524
rect 10928 17484 10934 17496
rect 11057 17493 11069 17496
rect 11103 17493 11115 17527
rect 11057 17487 11115 17493
rect 14093 17527 14151 17533
rect 14093 17493 14105 17527
rect 14139 17524 14151 17527
rect 15194 17524 15200 17536
rect 14139 17496 15200 17524
rect 14139 17493 14151 17496
rect 14093 17487 14151 17493
rect 15194 17484 15200 17496
rect 15252 17484 15258 17536
rect 18138 17484 18144 17536
rect 18196 17524 18202 17536
rect 18601 17527 18659 17533
rect 18601 17524 18613 17527
rect 18196 17496 18613 17524
rect 18196 17484 18202 17496
rect 18601 17493 18613 17496
rect 18647 17493 18659 17527
rect 18601 17487 18659 17493
rect 1104 17434 19136 17456
rect 1104 17382 3010 17434
rect 3062 17382 3074 17434
rect 3126 17382 3138 17434
rect 3190 17382 3202 17434
rect 3254 17382 3266 17434
rect 3318 17382 19136 17434
rect 1104 17360 19136 17382
rect 9214 17280 9220 17332
rect 9272 17320 9278 17332
rect 9309 17323 9367 17329
rect 9309 17320 9321 17323
rect 9272 17292 9321 17320
rect 9272 17280 9278 17292
rect 9309 17289 9321 17292
rect 9355 17289 9367 17323
rect 9309 17283 9367 17289
rect 10778 17280 10784 17332
rect 10836 17320 10842 17332
rect 11517 17323 11575 17329
rect 11517 17320 11529 17323
rect 10836 17292 11529 17320
rect 10836 17280 10842 17292
rect 11517 17289 11529 17292
rect 11563 17289 11575 17323
rect 11517 17283 11575 17289
rect 11882 17280 11888 17332
rect 11940 17280 11946 17332
rect 14737 17323 14795 17329
rect 14737 17289 14749 17323
rect 14783 17320 14795 17323
rect 14826 17320 14832 17332
rect 14783 17292 14832 17320
rect 14783 17289 14795 17292
rect 14737 17283 14795 17289
rect 14826 17280 14832 17292
rect 14884 17280 14890 17332
rect 15473 17323 15531 17329
rect 15473 17289 15485 17323
rect 15519 17320 15531 17323
rect 15746 17320 15752 17332
rect 15519 17292 15752 17320
rect 15519 17289 15531 17292
rect 15473 17283 15531 17289
rect 15746 17280 15752 17292
rect 15804 17280 15810 17332
rect 1210 17212 1216 17264
rect 1268 17252 1274 17264
rect 3421 17255 3479 17261
rect 3421 17252 3433 17255
rect 1268 17224 3433 17252
rect 1268 17212 1274 17224
rect 1578 17144 1584 17196
rect 1636 17144 1642 17196
rect 2130 17144 2136 17196
rect 2188 17184 2194 17196
rect 2314 17184 2320 17196
rect 2188 17156 2320 17184
rect 2188 17144 2194 17156
rect 2314 17144 2320 17156
rect 2372 17144 2378 17196
rect 2424 17193 2452 17224
rect 3421 17221 3433 17224
rect 3467 17221 3479 17255
rect 3421 17215 3479 17221
rect 6546 17212 6552 17264
rect 6604 17252 6610 17264
rect 7837 17255 7895 17261
rect 6604 17224 7604 17252
rect 6604 17212 6610 17224
rect 2409 17187 2467 17193
rect 2409 17153 2421 17187
rect 2455 17153 2467 17187
rect 2409 17147 2467 17153
rect 2501 17187 2559 17193
rect 2501 17153 2513 17187
rect 2547 17153 2559 17187
rect 2501 17147 2559 17153
rect 2685 17187 2743 17193
rect 2685 17153 2697 17187
rect 2731 17184 2743 17187
rect 2731 17156 3464 17184
rect 2731 17153 2743 17156
rect 2685 17147 2743 17153
rect 2222 17076 2228 17128
rect 2280 17116 2286 17128
rect 2516 17116 2544 17147
rect 2280 17088 2544 17116
rect 3436 17116 3464 17156
rect 3510 17144 3516 17196
rect 3568 17184 3574 17196
rect 4065 17187 4123 17193
rect 4065 17184 4077 17187
rect 3568 17156 4077 17184
rect 3568 17144 3574 17156
rect 4065 17153 4077 17156
rect 4111 17153 4123 17187
rect 4065 17147 4123 17153
rect 6181 17187 6239 17193
rect 6181 17153 6193 17187
rect 6227 17184 6239 17187
rect 6638 17184 6644 17196
rect 6227 17156 6644 17184
rect 6227 17153 6239 17156
rect 6181 17147 6239 17153
rect 6638 17144 6644 17156
rect 6696 17144 6702 17196
rect 7576 17193 7604 17224
rect 7837 17221 7849 17255
rect 7883 17252 7895 17255
rect 7926 17252 7932 17264
rect 7883 17224 7932 17252
rect 7883 17221 7895 17224
rect 7837 17215 7895 17221
rect 7926 17212 7932 17224
rect 7984 17212 7990 17264
rect 8570 17212 8576 17264
rect 8628 17212 8634 17264
rect 9858 17212 9864 17264
rect 9916 17212 9922 17264
rect 10870 17212 10876 17264
rect 10928 17212 10934 17264
rect 14918 17252 14924 17264
rect 12406 17224 14924 17252
rect 7561 17187 7619 17193
rect 7561 17153 7573 17187
rect 7607 17153 7619 17187
rect 7561 17147 7619 17153
rect 9582 17144 9588 17196
rect 9640 17144 9646 17196
rect 11422 17144 11428 17196
rect 11480 17184 11486 17196
rect 11517 17187 11575 17193
rect 11517 17184 11529 17187
rect 11480 17156 11529 17184
rect 11480 17144 11486 17156
rect 11517 17153 11529 17156
rect 11563 17153 11575 17187
rect 11517 17147 11575 17153
rect 11698 17144 11704 17196
rect 11756 17144 11762 17196
rect 12160 17187 12218 17193
rect 12160 17153 12172 17187
rect 12206 17153 12218 17187
rect 12160 17147 12218 17153
rect 3436 17088 3556 17116
rect 2280 17076 2286 17088
rect 3528 17060 3556 17088
rect 3878 17076 3884 17128
rect 3936 17076 3942 17128
rect 11330 17076 11336 17128
rect 11388 17076 11394 17128
rect 3510 17008 3516 17060
rect 3568 17008 3574 17060
rect 10962 17008 10968 17060
rect 11020 17048 11026 17060
rect 11716 17048 11744 17144
rect 12176 17116 12204 17147
rect 12250 17144 12256 17196
rect 12308 17184 12314 17196
rect 12406 17184 12434 17224
rect 14918 17212 14924 17224
rect 14976 17252 14982 17264
rect 18690 17252 18696 17264
rect 14976 17224 15148 17252
rect 14976 17212 14982 17224
rect 12308 17156 12434 17184
rect 12308 17144 12314 17156
rect 13722 17144 13728 17196
rect 13780 17184 13786 17196
rect 15120 17193 15148 17224
rect 17512 17224 18184 17252
rect 14829 17187 14887 17193
rect 14829 17184 14841 17187
rect 13780 17156 14841 17184
rect 13780 17144 13786 17156
rect 14829 17153 14841 17156
rect 14875 17153 14887 17187
rect 14829 17147 14887 17153
rect 15105 17187 15163 17193
rect 15105 17153 15117 17187
rect 15151 17153 15163 17187
rect 15105 17147 15163 17153
rect 15194 17144 15200 17196
rect 15252 17184 15258 17196
rect 15252 17156 15297 17184
rect 15252 17144 15258 17156
rect 17126 17144 17132 17196
rect 17184 17184 17190 17196
rect 17512 17193 17540 17224
rect 18156 17196 18184 17224
rect 18340 17224 18696 17252
rect 17497 17187 17555 17193
rect 17497 17184 17509 17187
rect 17184 17156 17509 17184
rect 17184 17144 17190 17156
rect 17497 17153 17509 17156
rect 17543 17153 17555 17187
rect 17497 17147 17555 17153
rect 17586 17144 17592 17196
rect 17644 17144 17650 17196
rect 17681 17187 17739 17193
rect 17681 17153 17693 17187
rect 17727 17153 17739 17187
rect 17681 17147 17739 17153
rect 12434 17116 12440 17128
rect 12176 17088 12440 17116
rect 12434 17076 12440 17088
rect 12492 17076 12498 17128
rect 17696 17116 17724 17147
rect 17770 17144 17776 17196
rect 17828 17184 17834 17196
rect 17865 17187 17923 17193
rect 17865 17184 17877 17187
rect 17828 17156 17877 17184
rect 17828 17144 17834 17156
rect 17865 17153 17877 17156
rect 17911 17153 17923 17187
rect 17865 17147 17923 17153
rect 18138 17144 18144 17196
rect 18196 17193 18202 17196
rect 18340 17193 18368 17224
rect 18690 17212 18696 17224
rect 18748 17212 18754 17264
rect 18196 17187 18229 17193
rect 18217 17153 18229 17187
rect 18196 17147 18229 17153
rect 18325 17187 18383 17193
rect 18325 17153 18337 17187
rect 18371 17153 18383 17187
rect 18325 17147 18383 17153
rect 18417 17187 18475 17193
rect 18417 17153 18429 17187
rect 18463 17153 18475 17187
rect 18417 17147 18475 17153
rect 18196 17144 18202 17147
rect 17957 17119 18015 17125
rect 17957 17116 17969 17119
rect 17696 17088 17969 17116
rect 17957 17085 17969 17088
rect 18003 17085 18015 17119
rect 18432 17116 18460 17147
rect 17957 17079 18015 17085
rect 18340 17088 18460 17116
rect 11020 17020 11744 17048
rect 11020 17008 11026 17020
rect 17862 17008 17868 17060
rect 17920 17048 17926 17060
rect 18340 17048 18368 17088
rect 17920 17020 18368 17048
rect 17920 17008 17926 17020
rect 1394 16940 1400 16992
rect 1452 16940 1458 16992
rect 2038 16940 2044 16992
rect 2096 16940 2102 16992
rect 2774 16940 2780 16992
rect 2832 16980 2838 16992
rect 3786 16980 3792 16992
rect 2832 16952 3792 16980
rect 2832 16940 2838 16952
rect 3786 16940 3792 16952
rect 3844 16940 3850 16992
rect 6086 16940 6092 16992
rect 6144 16940 6150 16992
rect 17221 16983 17279 16989
rect 17221 16949 17233 16983
rect 17267 16980 17279 16983
rect 17310 16980 17316 16992
rect 17267 16952 17316 16980
rect 17267 16949 17279 16952
rect 17221 16943 17279 16949
rect 17310 16940 17316 16952
rect 17368 16940 17374 16992
rect 18414 16940 18420 16992
rect 18472 16980 18478 16992
rect 18509 16983 18567 16989
rect 18509 16980 18521 16983
rect 18472 16952 18521 16980
rect 18472 16940 18478 16952
rect 18509 16949 18521 16952
rect 18555 16949 18567 16983
rect 18509 16943 18567 16949
rect 1104 16890 19136 16912
rect 1104 16838 2350 16890
rect 2402 16838 2414 16890
rect 2466 16838 2478 16890
rect 2530 16838 2542 16890
rect 2594 16838 2606 16890
rect 2658 16838 19136 16890
rect 1104 16816 19136 16838
rect 1397 16779 1455 16785
rect 1397 16745 1409 16779
rect 1443 16776 1455 16779
rect 1578 16776 1584 16788
rect 1443 16748 1584 16776
rect 1443 16745 1455 16748
rect 1397 16739 1455 16745
rect 1578 16736 1584 16748
rect 1636 16736 1642 16788
rect 1670 16736 1676 16788
rect 1728 16776 1734 16788
rect 1728 16748 4752 16776
rect 1728 16736 1734 16748
rect 3878 16668 3884 16720
rect 3936 16708 3942 16720
rect 4249 16711 4307 16717
rect 4249 16708 4261 16711
rect 3936 16680 4261 16708
rect 3936 16668 3942 16680
rect 4249 16677 4261 16680
rect 4295 16677 4307 16711
rect 4249 16671 4307 16677
rect 1670 16600 1676 16652
rect 1728 16600 1734 16652
rect 1949 16643 2007 16649
rect 1949 16609 1961 16643
rect 1995 16640 2007 16643
rect 2038 16640 2044 16652
rect 1995 16612 2044 16640
rect 1995 16609 2007 16612
rect 1949 16603 2007 16609
rect 2038 16600 2044 16612
rect 2096 16600 2102 16652
rect 3786 16600 3792 16652
rect 3844 16640 3850 16652
rect 4724 16649 4752 16748
rect 6454 16736 6460 16788
rect 6512 16736 6518 16788
rect 12618 16776 12624 16788
rect 10704 16748 12624 16776
rect 4709 16643 4767 16649
rect 3844 16612 4016 16640
rect 3844 16600 3850 16612
rect 1578 16532 1584 16584
rect 1636 16532 1642 16584
rect 3988 16581 4016 16612
rect 4709 16609 4721 16643
rect 4755 16609 4767 16643
rect 4709 16603 4767 16609
rect 4985 16643 5043 16649
rect 4985 16609 4997 16643
rect 5031 16640 5043 16643
rect 5718 16640 5724 16652
rect 5031 16612 5724 16640
rect 5031 16609 5043 16612
rect 4985 16603 5043 16609
rect 5718 16600 5724 16612
rect 5776 16600 5782 16652
rect 6546 16600 6552 16652
rect 6604 16600 6610 16652
rect 9582 16600 9588 16652
rect 9640 16640 9646 16652
rect 10704 16649 10732 16748
rect 12618 16736 12624 16748
rect 12676 16736 12682 16788
rect 12710 16736 12716 16788
rect 12768 16776 12774 16788
rect 13722 16776 13728 16788
rect 12768 16748 13728 16776
rect 12768 16736 12774 16748
rect 13722 16736 13728 16748
rect 13780 16776 13786 16788
rect 13780 16748 14504 16776
rect 13780 16736 13786 16748
rect 12406 16680 14136 16708
rect 10689 16643 10747 16649
rect 10689 16640 10701 16643
rect 9640 16612 10701 16640
rect 9640 16600 9646 16612
rect 10689 16609 10701 16612
rect 10735 16609 10747 16643
rect 10689 16603 10747 16609
rect 10962 16600 10968 16652
rect 11020 16600 11026 16652
rect 11422 16600 11428 16652
rect 11480 16640 11486 16652
rect 12406 16640 12434 16680
rect 11480 16612 12434 16640
rect 11480 16600 11486 16612
rect 3973 16575 4031 16581
rect 2774 16396 2780 16448
rect 2832 16436 2838 16448
rect 3068 16436 3096 16558
rect 3973 16541 3985 16575
rect 4019 16541 4031 16575
rect 3973 16535 4031 16541
rect 4524 16575 4582 16581
rect 4524 16541 4536 16575
rect 4570 16541 4582 16575
rect 4524 16535 4582 16541
rect 4540 16504 4568 16535
rect 4614 16532 4620 16584
rect 4672 16532 4678 16584
rect 6086 16532 6092 16584
rect 6144 16532 6150 16584
rect 6362 16532 6368 16584
rect 6420 16572 6426 16584
rect 8941 16575 8999 16581
rect 8941 16572 8953 16575
rect 6420 16544 8953 16572
rect 6420 16532 6426 16544
rect 8941 16541 8953 16544
rect 8987 16541 8999 16575
rect 8941 16535 8999 16541
rect 9095 16575 9153 16581
rect 9095 16541 9107 16575
rect 9141 16572 9153 16575
rect 9214 16572 9220 16584
rect 9141 16544 9220 16572
rect 9141 16541 9153 16544
rect 9095 16535 9153 16541
rect 4890 16504 4896 16516
rect 4540 16476 4896 16504
rect 4890 16464 4896 16476
rect 4948 16464 4954 16516
rect 8294 16464 8300 16516
rect 8352 16464 8358 16516
rect 8956 16504 8984 16535
rect 9214 16532 9220 16544
rect 9272 16532 9278 16584
rect 12710 16532 12716 16584
rect 12768 16532 12774 16584
rect 14108 16581 14136 16680
rect 14476 16581 14504 16748
rect 18690 16736 18696 16788
rect 18748 16776 18754 16788
rect 18785 16779 18843 16785
rect 18785 16776 18797 16779
rect 18748 16748 18797 16776
rect 18748 16736 18754 16748
rect 18785 16745 18797 16748
rect 18831 16745 18843 16779
rect 18785 16739 18843 16745
rect 15838 16600 15844 16652
rect 15896 16640 15902 16652
rect 17037 16643 17095 16649
rect 17037 16640 17049 16643
rect 15896 16612 17049 16640
rect 15896 16600 15902 16612
rect 17037 16609 17049 16612
rect 17083 16609 17095 16643
rect 17037 16603 17095 16609
rect 17310 16600 17316 16652
rect 17368 16600 17374 16652
rect 14093 16575 14151 16581
rect 14093 16541 14105 16575
rect 14139 16541 14151 16575
rect 14093 16535 14151 16541
rect 14277 16575 14335 16581
rect 14277 16541 14289 16575
rect 14323 16541 14335 16575
rect 14277 16535 14335 16541
rect 14461 16575 14519 16581
rect 14461 16541 14473 16575
rect 14507 16541 14519 16575
rect 14461 16535 14519 16541
rect 12621 16507 12679 16513
rect 12621 16504 12633 16507
rect 8956 16476 11376 16504
rect 12190 16476 12633 16504
rect 2832 16408 3096 16436
rect 2832 16396 2838 16408
rect 3418 16396 3424 16448
rect 3476 16396 3482 16448
rect 4062 16396 4068 16448
rect 4120 16396 4126 16448
rect 4614 16396 4620 16448
rect 4672 16436 4678 16448
rect 6362 16436 6368 16448
rect 4672 16408 6368 16436
rect 4672 16396 4678 16408
rect 6362 16396 6368 16408
rect 6420 16396 6426 16448
rect 6638 16396 6644 16448
rect 6696 16436 6702 16448
rect 8662 16436 8668 16448
rect 6696 16408 8668 16436
rect 6696 16396 6702 16408
rect 8662 16396 8668 16408
rect 8720 16396 8726 16448
rect 9309 16439 9367 16445
rect 9309 16405 9321 16439
rect 9355 16436 9367 16439
rect 9490 16436 9496 16448
rect 9355 16408 9496 16436
rect 9355 16405 9367 16408
rect 9309 16399 9367 16405
rect 9490 16396 9496 16408
rect 9548 16396 9554 16448
rect 11348 16436 11376 16476
rect 12621 16473 12633 16476
rect 12667 16473 12679 16507
rect 14292 16504 14320 16535
rect 14918 16532 14924 16584
rect 14976 16532 14982 16584
rect 15010 16532 15016 16584
rect 15068 16532 15074 16584
rect 18414 16532 18420 16584
rect 18472 16532 18478 16584
rect 14292 16476 17172 16504
rect 12621 16467 12679 16473
rect 17144 16448 17172 16476
rect 12250 16436 12256 16448
rect 11348 16408 12256 16436
rect 12250 16396 12256 16408
rect 12308 16396 12314 16448
rect 12434 16396 12440 16448
rect 12492 16396 12498 16448
rect 14185 16439 14243 16445
rect 14185 16405 14197 16439
rect 14231 16436 14243 16439
rect 14458 16436 14464 16448
rect 14231 16408 14464 16436
rect 14231 16405 14243 16408
rect 14185 16399 14243 16405
rect 14458 16396 14464 16408
rect 14516 16396 14522 16448
rect 14550 16396 14556 16448
rect 14608 16396 14614 16448
rect 15289 16439 15347 16445
rect 15289 16405 15301 16439
rect 15335 16436 15347 16439
rect 16206 16436 16212 16448
rect 15335 16408 16212 16436
rect 15335 16405 15347 16408
rect 15289 16399 15347 16405
rect 16206 16396 16212 16408
rect 16264 16396 16270 16448
rect 17126 16396 17132 16448
rect 17184 16396 17190 16448
rect 1104 16346 19136 16368
rect 1104 16294 3010 16346
rect 3062 16294 3074 16346
rect 3126 16294 3138 16346
rect 3190 16294 3202 16346
rect 3254 16294 3266 16346
rect 3318 16294 19136 16346
rect 1104 16272 19136 16294
rect 2222 16192 2228 16244
rect 2280 16232 2286 16244
rect 2409 16235 2467 16241
rect 2409 16232 2421 16235
rect 2280 16204 2421 16232
rect 2280 16192 2286 16204
rect 2409 16201 2421 16204
rect 2455 16201 2467 16235
rect 2409 16195 2467 16201
rect 2774 16192 2780 16244
rect 2832 16192 2838 16244
rect 4890 16192 4896 16244
rect 4948 16192 4954 16244
rect 8386 16232 8392 16244
rect 7760 16204 8392 16232
rect 1578 16124 1584 16176
rect 1636 16164 1642 16176
rect 3418 16164 3424 16176
rect 1636 16136 3424 16164
rect 1636 16124 1642 16136
rect 842 16056 848 16108
rect 900 16096 906 16108
rect 2056 16105 2084 16136
rect 3418 16124 3424 16136
rect 3476 16124 3482 16176
rect 4062 16124 4068 16176
rect 4120 16124 4126 16176
rect 7760 16173 7788 16204
rect 8386 16192 8392 16204
rect 8444 16192 8450 16244
rect 9214 16192 9220 16244
rect 9272 16192 9278 16244
rect 12618 16192 12624 16244
rect 12676 16232 12682 16244
rect 15473 16235 15531 16241
rect 15473 16232 15485 16235
rect 12676 16204 15485 16232
rect 12676 16192 12682 16204
rect 15473 16201 15485 16204
rect 15519 16232 15531 16235
rect 15838 16232 15844 16244
rect 15519 16204 15844 16232
rect 15519 16201 15531 16204
rect 15473 16195 15531 16201
rect 15838 16192 15844 16204
rect 15896 16192 15902 16244
rect 18417 16235 18475 16241
rect 18417 16201 18429 16235
rect 18463 16232 18475 16235
rect 18506 16232 18512 16244
rect 18463 16204 18512 16232
rect 18463 16201 18475 16204
rect 18417 16195 18475 16201
rect 18506 16192 18512 16204
rect 18564 16192 18570 16244
rect 7745 16167 7803 16173
rect 7745 16164 7757 16167
rect 7208 16136 7757 16164
rect 1397 16099 1455 16105
rect 1397 16096 1409 16099
rect 900 16068 1409 16096
rect 900 16056 906 16068
rect 1397 16065 1409 16068
rect 1443 16065 1455 16099
rect 1397 16059 1455 16065
rect 2041 16099 2099 16105
rect 2041 16065 2053 16099
rect 2087 16065 2099 16099
rect 2041 16059 2099 16065
rect 2130 16056 2136 16108
rect 2188 16056 2194 16108
rect 2682 16056 2688 16108
rect 2740 16056 2746 16108
rect 2866 16056 2872 16108
rect 2924 16096 2930 16108
rect 3145 16099 3203 16105
rect 3145 16096 3157 16099
rect 2924 16068 3157 16096
rect 2924 16056 2930 16068
rect 3145 16065 3157 16068
rect 3191 16065 3203 16099
rect 3145 16059 3203 16065
rect 6914 16056 6920 16108
rect 6972 16096 6978 16108
rect 7208 16105 7236 16136
rect 7745 16133 7757 16136
rect 7791 16133 7803 16167
rect 7745 16127 7803 16133
rect 8478 16124 8484 16176
rect 8536 16124 8542 16176
rect 13262 16124 13268 16176
rect 13320 16124 13326 16176
rect 17494 16124 17500 16176
rect 17552 16124 17558 16176
rect 7193 16099 7251 16105
rect 7193 16096 7205 16099
rect 6972 16068 7205 16096
rect 6972 16056 6978 16068
rect 7193 16065 7205 16068
rect 7239 16065 7251 16099
rect 7193 16059 7251 16065
rect 7374 16056 7380 16108
rect 7432 16056 7438 16108
rect 9490 16056 9496 16108
rect 9548 16056 9554 16108
rect 14182 16056 14188 16108
rect 14240 16056 14246 16108
rect 15930 16056 15936 16108
rect 15988 16096 15994 16108
rect 16669 16099 16727 16105
rect 16669 16096 16681 16099
rect 15988 16068 16681 16096
rect 15988 16056 15994 16068
rect 16669 16065 16681 16068
rect 16715 16065 16727 16099
rect 16669 16059 16727 16065
rect 18782 16056 18788 16108
rect 18840 16056 18846 16108
rect 2148 15960 2176 16056
rect 3421 16031 3479 16037
rect 3421 16028 3433 16031
rect 2746 16000 3433 16028
rect 2746 15960 2774 16000
rect 3421 15997 3433 16000
rect 3467 15997 3479 16031
rect 3421 15991 3479 15997
rect 6546 15988 6552 16040
rect 6604 16028 6610 16040
rect 7469 16031 7527 16037
rect 7469 16028 7481 16031
rect 6604 16000 7481 16028
rect 6604 15988 6610 16000
rect 7469 15997 7481 16000
rect 7515 15997 7527 16031
rect 7469 15991 7527 15997
rect 8110 15988 8116 16040
rect 8168 16028 8174 16040
rect 9309 16031 9367 16037
rect 9309 16028 9321 16031
rect 8168 16000 9321 16028
rect 8168 15988 8174 16000
rect 9309 15997 9321 16000
rect 9355 15997 9367 16031
rect 9309 15991 9367 15997
rect 12345 16031 12403 16037
rect 12345 15997 12357 16031
rect 12391 15997 12403 16031
rect 12345 15991 12403 15997
rect 12621 16031 12679 16037
rect 12621 15997 12633 16031
rect 12667 16028 12679 16031
rect 14090 16028 14096 16040
rect 12667 16000 14096 16028
rect 12667 15997 12679 16000
rect 12621 15991 12679 15997
rect 2148 15932 2774 15960
rect 9674 15920 9680 15972
rect 9732 15920 9738 15972
rect 1581 15895 1639 15901
rect 1581 15861 1593 15895
rect 1627 15892 1639 15895
rect 1762 15892 1768 15904
rect 1627 15864 1768 15892
rect 1627 15861 1639 15864
rect 1581 15855 1639 15861
rect 1762 15852 1768 15864
rect 1820 15852 1826 15904
rect 2682 15852 2688 15904
rect 2740 15892 2746 15904
rect 5810 15892 5816 15904
rect 2740 15864 5816 15892
rect 2740 15852 2746 15864
rect 5810 15852 5816 15864
rect 5868 15852 5874 15904
rect 7282 15852 7288 15904
rect 7340 15852 7346 15904
rect 12360 15892 12388 15991
rect 14090 15988 14096 16000
rect 14148 15988 14154 16040
rect 16945 16031 17003 16037
rect 16945 15997 16957 16031
rect 16991 16028 17003 16031
rect 17310 16028 17316 16040
rect 16991 16000 17316 16028
rect 16991 15997 17003 16000
rect 16945 15991 17003 15997
rect 17310 15988 17316 16000
rect 17368 15988 17374 16040
rect 13354 15892 13360 15904
rect 12360 15864 13360 15892
rect 13354 15852 13360 15864
rect 13412 15852 13418 15904
rect 14093 15895 14151 15901
rect 14093 15861 14105 15895
rect 14139 15892 14151 15895
rect 14366 15892 14372 15904
rect 14139 15864 14372 15892
rect 14139 15861 14151 15864
rect 14093 15855 14151 15861
rect 14366 15852 14372 15864
rect 14424 15852 14430 15904
rect 18138 15852 18144 15904
rect 18196 15892 18202 15904
rect 18601 15895 18659 15901
rect 18601 15892 18613 15895
rect 18196 15864 18613 15892
rect 18196 15852 18202 15864
rect 18601 15861 18613 15864
rect 18647 15861 18659 15895
rect 18601 15855 18659 15861
rect 1104 15802 19136 15824
rect 1104 15750 2350 15802
rect 2402 15750 2414 15802
rect 2466 15750 2478 15802
rect 2530 15750 2542 15802
rect 2594 15750 2606 15802
rect 2658 15750 19136 15802
rect 1104 15728 19136 15750
rect 6638 15688 6644 15700
rect 6196 15660 6644 15688
rect 2317 15623 2375 15629
rect 2317 15589 2329 15623
rect 2363 15589 2375 15623
rect 2317 15583 2375 15589
rect 1581 15487 1639 15493
rect 1581 15453 1593 15487
rect 1627 15484 1639 15487
rect 2332 15484 2360 15583
rect 1627 15456 2360 15484
rect 2501 15487 2559 15493
rect 1627 15453 1639 15456
rect 1581 15447 1639 15453
rect 2501 15453 2513 15487
rect 2547 15484 2559 15487
rect 3418 15484 3424 15496
rect 2547 15456 3424 15484
rect 2547 15453 2559 15456
rect 2501 15447 2559 15453
rect 3418 15444 3424 15456
rect 3476 15444 3482 15496
rect 5810 15444 5816 15496
rect 5868 15484 5874 15496
rect 6196 15484 6224 15660
rect 6638 15648 6644 15660
rect 6696 15648 6702 15700
rect 8021 15691 8079 15697
rect 8021 15657 8033 15691
rect 8067 15688 8079 15691
rect 8110 15688 8116 15700
rect 8067 15660 8116 15688
rect 8067 15657 8079 15660
rect 8021 15651 8079 15657
rect 8110 15648 8116 15660
rect 8168 15648 8174 15700
rect 8478 15648 8484 15700
rect 8536 15688 8542 15700
rect 8573 15691 8631 15697
rect 8573 15688 8585 15691
rect 8536 15660 8585 15688
rect 8536 15648 8542 15660
rect 8573 15657 8585 15660
rect 8619 15657 8631 15691
rect 8573 15651 8631 15657
rect 10781 15691 10839 15697
rect 10781 15657 10793 15691
rect 10827 15688 10839 15691
rect 11514 15688 11520 15700
rect 10827 15660 11520 15688
rect 10827 15657 10839 15660
rect 10781 15651 10839 15657
rect 11514 15648 11520 15660
rect 11572 15648 11578 15700
rect 13262 15648 13268 15700
rect 13320 15688 13326 15700
rect 13357 15691 13415 15697
rect 13357 15688 13369 15691
rect 13320 15660 13369 15688
rect 13320 15648 13326 15660
rect 13357 15657 13369 15660
rect 13403 15657 13415 15691
rect 13357 15651 13415 15657
rect 14185 15691 14243 15697
rect 14185 15657 14197 15691
rect 14231 15688 14243 15691
rect 15010 15688 15016 15700
rect 14231 15660 15016 15688
rect 14231 15657 14243 15660
rect 14185 15651 14243 15657
rect 15010 15648 15016 15660
rect 15068 15648 15074 15700
rect 17126 15688 17132 15700
rect 16592 15660 17132 15688
rect 16592 15620 16620 15660
rect 17126 15648 17132 15660
rect 17184 15648 17190 15700
rect 17494 15648 17500 15700
rect 17552 15648 17558 15700
rect 15856 15592 16620 15620
rect 16669 15623 16727 15629
rect 6273 15555 6331 15561
rect 6273 15521 6285 15555
rect 6319 15552 6331 15555
rect 6546 15552 6552 15564
rect 6319 15524 6552 15552
rect 6319 15521 6331 15524
rect 6273 15515 6331 15521
rect 6546 15512 6552 15524
rect 6604 15552 6610 15564
rect 9033 15555 9091 15561
rect 9033 15552 9045 15555
rect 6604 15524 9045 15552
rect 6604 15512 6610 15524
rect 9033 15521 9045 15524
rect 9079 15521 9091 15555
rect 12710 15552 12716 15564
rect 9033 15515 9091 15521
rect 12406 15524 12716 15552
rect 5868 15456 6224 15484
rect 8297 15487 8355 15493
rect 5868 15444 5874 15456
rect 8297 15453 8309 15487
rect 8343 15484 8355 15487
rect 8481 15487 8539 15493
rect 8481 15484 8493 15487
rect 8343 15456 8493 15484
rect 8343 15453 8355 15456
rect 8297 15447 8355 15453
rect 8481 15453 8493 15456
rect 8527 15453 8539 15487
rect 8481 15447 8539 15453
rect 11057 15487 11115 15493
rect 11057 15453 11069 15487
rect 11103 15484 11115 15487
rect 12406 15484 12434 15524
rect 12710 15512 12716 15524
rect 12768 15552 12774 15564
rect 15657 15555 15715 15561
rect 12768 15524 13308 15552
rect 12768 15512 12774 15524
rect 11103 15456 12434 15484
rect 11103 15453 11115 15456
rect 11057 15447 11115 15453
rect 6549 15419 6607 15425
rect 6549 15385 6561 15419
rect 6595 15385 6607 15419
rect 8205 15419 8263 15425
rect 8205 15416 8217 15419
rect 7774 15388 8217 15416
rect 6549 15379 6607 15385
rect 8205 15385 8217 15388
rect 8251 15385 8263 15419
rect 8205 15379 8263 15385
rect 1394 15308 1400 15360
rect 1452 15308 1458 15360
rect 2130 15308 2136 15360
rect 2188 15348 2194 15360
rect 2682 15348 2688 15360
rect 2188 15320 2688 15348
rect 2188 15308 2194 15320
rect 2682 15308 2688 15320
rect 2740 15308 2746 15360
rect 5718 15308 5724 15360
rect 5776 15308 5782 15360
rect 6564 15348 6592 15379
rect 7190 15348 7196 15360
rect 6564 15320 7196 15348
rect 7190 15308 7196 15320
rect 7248 15308 7254 15360
rect 8496 15348 8524 15447
rect 9306 15376 9312 15428
rect 9364 15376 9370 15428
rect 10965 15419 11023 15425
rect 10965 15416 10977 15419
rect 10534 15388 10977 15416
rect 10965 15385 10977 15388
rect 11011 15385 11023 15419
rect 10965 15379 11023 15385
rect 8662 15348 8668 15360
rect 8496 15320 8668 15348
rect 8662 15308 8668 15320
rect 8720 15348 8726 15360
rect 11072 15348 11100 15447
rect 12618 15444 12624 15496
rect 12676 15484 12682 15496
rect 13280 15493 13308 15524
rect 15657 15521 15669 15555
rect 15703 15552 15715 15555
rect 15856 15552 15884 15592
rect 16669 15589 16681 15623
rect 16715 15620 16727 15623
rect 17586 15620 17592 15632
rect 16715 15592 17592 15620
rect 16715 15589 16727 15592
rect 16669 15583 16727 15589
rect 17586 15580 17592 15592
rect 17644 15580 17650 15632
rect 15703 15524 15884 15552
rect 15703 15521 15715 15524
rect 15657 15515 15715 15521
rect 15930 15512 15936 15564
rect 15988 15512 15994 15564
rect 16206 15512 16212 15564
rect 16264 15512 16270 15564
rect 12989 15487 13047 15493
rect 12989 15484 13001 15487
rect 12676 15456 13001 15484
rect 12676 15444 12682 15456
rect 12989 15453 13001 15456
rect 13035 15453 13047 15487
rect 12989 15447 13047 15453
rect 13265 15487 13323 15493
rect 13265 15453 13277 15487
rect 13311 15484 13323 15487
rect 13722 15484 13728 15496
rect 13311 15456 13728 15484
rect 13311 15453 13323 15456
rect 13265 15447 13323 15453
rect 13722 15444 13728 15456
rect 13780 15444 13786 15496
rect 14550 15444 14556 15496
rect 14608 15444 14614 15496
rect 16025 15487 16083 15493
rect 16025 15484 16037 15487
rect 15948 15456 16037 15484
rect 8720 15320 11100 15348
rect 8720 15308 8726 15320
rect 14366 15308 14372 15360
rect 14424 15348 14430 15360
rect 15948 15348 15976 15456
rect 16025 15453 16037 15456
rect 16071 15453 16083 15487
rect 16025 15447 16083 15453
rect 16758 15444 16764 15496
rect 16816 15444 16822 15496
rect 17405 15487 17463 15493
rect 17405 15453 17417 15487
rect 17451 15484 17463 15487
rect 17494 15484 17500 15496
rect 17451 15456 17500 15484
rect 17451 15453 17463 15456
rect 17405 15447 17463 15453
rect 17494 15444 17500 15456
rect 17552 15484 17558 15496
rect 17862 15484 17868 15496
rect 17552 15456 17868 15484
rect 17552 15444 17558 15456
rect 17862 15444 17868 15456
rect 17920 15444 17926 15496
rect 18322 15444 18328 15496
rect 18380 15484 18386 15496
rect 18601 15487 18659 15493
rect 18601 15484 18613 15487
rect 18380 15456 18613 15484
rect 18380 15444 18386 15456
rect 18601 15453 18613 15456
rect 18647 15453 18659 15487
rect 18601 15447 18659 15453
rect 17129 15419 17187 15425
rect 17129 15385 17141 15419
rect 17175 15416 17187 15419
rect 18506 15416 18512 15428
rect 17175 15388 18512 15416
rect 17175 15385 17187 15388
rect 17129 15379 17187 15385
rect 18506 15376 18512 15388
rect 18564 15376 18570 15428
rect 14424 15320 15976 15348
rect 14424 15308 14430 15320
rect 17310 15308 17316 15360
rect 17368 15308 17374 15360
rect 18782 15308 18788 15360
rect 18840 15308 18846 15360
rect 1104 15258 19136 15280
rect 1104 15206 3010 15258
rect 3062 15206 3074 15258
rect 3126 15206 3138 15258
rect 3190 15206 3202 15258
rect 3254 15206 3266 15258
rect 3318 15206 19136 15258
rect 1104 15184 19136 15206
rect 1854 15144 1860 15156
rect 1412 15116 1860 15144
rect 1412 15017 1440 15116
rect 1854 15104 1860 15116
rect 1912 15144 1918 15156
rect 3145 15147 3203 15153
rect 1912 15116 3004 15144
rect 1912 15104 1918 15116
rect 2976 15088 3004 15116
rect 3145 15113 3157 15147
rect 3191 15144 3203 15147
rect 3418 15144 3424 15156
rect 3191 15116 3424 15144
rect 3191 15113 3203 15116
rect 3145 15107 3203 15113
rect 3418 15104 3424 15116
rect 3476 15104 3482 15156
rect 7101 15147 7159 15153
rect 7101 15113 7113 15147
rect 7147 15113 7159 15147
rect 7101 15107 7159 15113
rect 2958 15036 2964 15088
rect 3016 15076 3022 15088
rect 5718 15076 5724 15088
rect 3016 15048 3832 15076
rect 5290 15048 5724 15076
rect 3016 15036 3022 15048
rect 3804 15020 3832 15048
rect 5718 15036 5724 15048
rect 5776 15036 5782 15088
rect 6917 15079 6975 15085
rect 6917 15045 6929 15079
rect 6963 15076 6975 15079
rect 7006 15076 7012 15088
rect 6963 15048 7012 15076
rect 6963 15045 6975 15048
rect 6917 15039 6975 15045
rect 7006 15036 7012 15048
rect 7064 15036 7070 15088
rect 7116 15076 7144 15107
rect 7190 15104 7196 15156
rect 7248 15104 7254 15156
rect 7282 15104 7288 15156
rect 7340 15144 7346 15156
rect 7561 15147 7619 15153
rect 7561 15144 7573 15147
rect 7340 15116 7573 15144
rect 7340 15104 7346 15116
rect 7561 15113 7573 15116
rect 7607 15113 7619 15147
rect 7561 15107 7619 15113
rect 14090 15104 14096 15156
rect 14148 15104 14154 15156
rect 14458 15104 14464 15156
rect 14516 15104 14522 15156
rect 9306 15076 9312 15088
rect 7116 15048 9312 15076
rect 1397 15011 1455 15017
rect 1397 14977 1409 15011
rect 1443 14977 1455 15011
rect 1397 14971 1455 14977
rect 2774 14968 2780 15020
rect 2832 14968 2838 15020
rect 3513 15011 3571 15017
rect 3513 15008 3525 15011
rect 2884 14980 3525 15008
rect 1670 14900 1676 14952
rect 1728 14900 1734 14952
rect 1762 14900 1768 14952
rect 1820 14940 1826 14952
rect 2682 14940 2688 14952
rect 1820 14912 2688 14940
rect 1820 14900 1826 14912
rect 2682 14900 2688 14912
rect 2740 14940 2746 14952
rect 2884 14940 2912 14980
rect 3513 14977 3525 14980
rect 3559 14977 3571 15011
rect 3513 14971 3571 14977
rect 3694 14968 3700 15020
rect 3752 14968 3758 15020
rect 3786 14968 3792 15020
rect 3844 14968 3850 15020
rect 5626 14968 5632 15020
rect 5684 14968 5690 15020
rect 7392 15017 7420 15048
rect 9306 15036 9312 15048
rect 9364 15036 9370 15088
rect 11422 15036 11428 15088
rect 11480 15076 11486 15088
rect 11701 15079 11759 15085
rect 11701 15076 11713 15079
rect 11480 15048 11713 15076
rect 11480 15036 11486 15048
rect 11701 15045 11713 15048
rect 11747 15045 11759 15079
rect 17310 15076 17316 15088
rect 11701 15039 11759 15045
rect 14292 15048 17316 15076
rect 7377 15011 7435 15017
rect 7377 14977 7389 15011
rect 7423 14977 7435 15011
rect 7377 14971 7435 14977
rect 7653 15011 7711 15017
rect 7653 14977 7665 15011
rect 7699 15008 7711 15011
rect 8110 15008 8116 15020
rect 7699 14980 8116 15008
rect 7699 14977 7711 14980
rect 7653 14971 7711 14977
rect 8110 14968 8116 14980
rect 8168 14968 8174 15020
rect 11790 14968 11796 15020
rect 11848 14968 11854 15020
rect 14292 15017 14320 15048
rect 17310 15036 17316 15048
rect 17368 15036 17374 15088
rect 17420 15048 17908 15076
rect 14277 15011 14335 15017
rect 14277 14977 14289 15011
rect 14323 14977 14335 15011
rect 14277 14971 14335 14977
rect 14366 14968 14372 15020
rect 14424 15008 14430 15020
rect 14553 15011 14611 15017
rect 14553 15008 14565 15011
rect 14424 14980 14565 15008
rect 14424 14968 14430 14980
rect 14553 14977 14565 14980
rect 14599 14977 14611 15011
rect 14553 14971 14611 14977
rect 17034 14968 17040 15020
rect 17092 15008 17098 15020
rect 17420 15017 17448 15048
rect 17405 15011 17463 15017
rect 17405 15008 17417 15011
rect 17092 14980 17417 15008
rect 17092 14968 17098 14980
rect 17405 14977 17417 14980
rect 17451 14977 17463 15011
rect 17405 14971 17463 14977
rect 17497 15011 17555 15017
rect 17497 14977 17509 15011
rect 17543 14977 17555 15011
rect 17497 14971 17555 14977
rect 17589 15011 17647 15017
rect 17589 14977 17601 15011
rect 17635 14977 17647 15011
rect 17589 14971 17647 14977
rect 2740 14912 2912 14940
rect 2740 14900 2746 14912
rect 4062 14900 4068 14952
rect 4120 14900 4126 14952
rect 4522 14900 4528 14952
rect 4580 14940 4586 14952
rect 6549 14943 6607 14949
rect 6549 14940 6561 14943
rect 4580 14912 6561 14940
rect 4580 14900 4586 14912
rect 6549 14909 6561 14912
rect 6595 14940 6607 14943
rect 11808 14940 11836 14968
rect 6595 14912 11836 14940
rect 6595 14909 6607 14912
rect 6549 14903 6607 14909
rect 15470 14900 15476 14952
rect 15528 14900 15534 14952
rect 15654 14900 15660 14952
rect 15712 14900 15718 14952
rect 16117 14943 16175 14949
rect 16117 14909 16129 14943
rect 16163 14940 16175 14943
rect 17512 14940 17540 14971
rect 16163 14912 17540 14940
rect 17604 14940 17632 14971
rect 17770 14968 17776 15020
rect 17828 14968 17834 15020
rect 17880 15008 17908 15048
rect 18138 15008 18144 15020
rect 17880 14980 18144 15008
rect 18138 14968 18144 14980
rect 18196 14968 18202 15020
rect 18230 14968 18236 15020
rect 18288 14968 18294 15020
rect 18785 15011 18843 15017
rect 18785 14977 18797 15011
rect 18831 15008 18843 15011
rect 18874 15008 18880 15020
rect 18831 14980 18880 15008
rect 18831 14977 18843 14980
rect 18785 14971 18843 14977
rect 18874 14968 18880 14980
rect 18932 14968 18938 15020
rect 17865 14943 17923 14949
rect 17865 14940 17877 14943
rect 17604 14912 17877 14940
rect 16163 14909 16175 14912
rect 16117 14903 16175 14909
rect 17512 14872 17540 14912
rect 17865 14909 17877 14912
rect 17911 14909 17923 14943
rect 17865 14903 17923 14909
rect 17954 14872 17960 14884
rect 17512 14844 17960 14872
rect 17954 14832 17960 14844
rect 18012 14832 18018 14884
rect 3602 14764 3608 14816
rect 3660 14764 3666 14816
rect 5534 14764 5540 14816
rect 5592 14764 5598 14816
rect 6914 14764 6920 14816
rect 6972 14764 6978 14816
rect 17129 14807 17187 14813
rect 17129 14773 17141 14807
rect 17175 14804 17187 14807
rect 17310 14804 17316 14816
rect 17175 14776 17316 14804
rect 17175 14773 17187 14776
rect 17129 14767 17187 14773
rect 17310 14764 17316 14776
rect 17368 14764 17374 14816
rect 17402 14764 17408 14816
rect 17460 14804 17466 14816
rect 18601 14807 18659 14813
rect 18601 14804 18613 14807
rect 17460 14776 18613 14804
rect 17460 14764 17466 14776
rect 18601 14773 18613 14776
rect 18647 14773 18659 14807
rect 18601 14767 18659 14773
rect 1104 14714 19136 14736
rect 1104 14662 2350 14714
rect 2402 14662 2414 14714
rect 2466 14662 2478 14714
rect 2530 14662 2542 14714
rect 2594 14662 2606 14714
rect 2658 14662 19136 14714
rect 1104 14640 19136 14662
rect 2501 14603 2559 14609
rect 2501 14569 2513 14603
rect 2547 14600 2559 14603
rect 2774 14600 2780 14612
rect 2547 14572 2780 14600
rect 2547 14569 2559 14572
rect 2501 14563 2559 14569
rect 2774 14560 2780 14572
rect 2832 14560 2838 14612
rect 3789 14603 3847 14609
rect 3789 14569 3801 14603
rect 3835 14600 3847 14603
rect 4062 14600 4068 14612
rect 3835 14572 4068 14600
rect 3835 14569 3847 14572
rect 3789 14563 3847 14569
rect 4062 14560 4068 14572
rect 4120 14560 4126 14612
rect 14642 14560 14648 14612
rect 14700 14600 14706 14612
rect 14700 14572 14872 14600
rect 14700 14560 14706 14572
rect 1946 14492 1952 14544
rect 2004 14532 2010 14544
rect 2225 14535 2283 14541
rect 2225 14532 2237 14535
rect 2004 14504 2237 14532
rect 2004 14492 2010 14504
rect 2225 14501 2237 14504
rect 2271 14532 2283 14535
rect 3510 14532 3516 14544
rect 2271 14504 3516 14532
rect 2271 14501 2283 14504
rect 2225 14495 2283 14501
rect 3510 14492 3516 14504
rect 3568 14492 3574 14544
rect 3694 14492 3700 14544
rect 3752 14532 3758 14544
rect 4341 14535 4399 14541
rect 4341 14532 4353 14535
rect 3752 14504 4353 14532
rect 3752 14492 3758 14504
rect 4341 14501 4353 14504
rect 4387 14501 4399 14535
rect 4341 14495 4399 14501
rect 13354 14492 13360 14544
rect 13412 14532 13418 14544
rect 13412 14504 14780 14532
rect 13412 14492 13418 14504
rect 1489 14467 1547 14473
rect 1489 14433 1501 14467
rect 1535 14464 1547 14467
rect 1670 14464 1676 14476
rect 1535 14436 1676 14464
rect 1535 14433 1547 14436
rect 1489 14427 1547 14433
rect 1670 14424 1676 14436
rect 1728 14464 1734 14476
rect 1728 14436 2774 14464
rect 1728 14424 1734 14436
rect 1762 14356 1768 14408
rect 1820 14356 1826 14408
rect 2130 14356 2136 14408
rect 2188 14396 2194 14408
rect 2409 14399 2467 14405
rect 2409 14396 2421 14399
rect 2188 14368 2421 14396
rect 2188 14356 2194 14368
rect 2409 14365 2421 14368
rect 2455 14365 2467 14399
rect 2746 14396 2774 14436
rect 3786 14424 3792 14476
rect 3844 14464 3850 14476
rect 5077 14467 5135 14473
rect 5077 14464 5089 14467
rect 3844 14436 5089 14464
rect 3844 14424 3850 14436
rect 5077 14433 5089 14436
rect 5123 14464 5135 14467
rect 5626 14464 5632 14476
rect 5123 14436 5632 14464
rect 5123 14433 5135 14436
rect 5077 14427 5135 14433
rect 5626 14424 5632 14436
rect 5684 14424 5690 14476
rect 11422 14424 11428 14476
rect 11480 14464 11486 14476
rect 14752 14473 14780 14504
rect 14744 14467 14802 14473
rect 11480 14436 14504 14464
rect 11480 14424 11486 14436
rect 3973 14399 4031 14405
rect 3973 14396 3985 14399
rect 2746 14368 3985 14396
rect 2409 14359 2467 14365
rect 3973 14365 3985 14368
rect 4019 14365 4031 14399
rect 3973 14359 4031 14365
rect 4249 14399 4307 14405
rect 4249 14365 4261 14399
rect 4295 14365 4307 14399
rect 4249 14359 4307 14365
rect 2225 14331 2283 14337
rect 2225 14328 2237 14331
rect 1780 14300 2237 14328
rect 1780 14272 1808 14300
rect 2225 14297 2237 14300
rect 2271 14297 2283 14331
rect 2225 14291 2283 14297
rect 3602 14288 3608 14340
rect 3660 14328 3666 14340
rect 4157 14331 4215 14337
rect 4157 14328 4169 14331
rect 3660 14300 4169 14328
rect 3660 14288 3666 14300
rect 4157 14297 4169 14300
rect 4203 14297 4215 14331
rect 4264 14328 4292 14359
rect 4338 14356 4344 14408
rect 4396 14356 4402 14408
rect 4522 14356 4528 14408
rect 4580 14356 4586 14408
rect 6825 14399 6883 14405
rect 6825 14365 6837 14399
rect 6871 14396 6883 14399
rect 8294 14396 8300 14408
rect 6871 14368 8300 14396
rect 6871 14365 6883 14368
rect 6825 14359 6883 14365
rect 8294 14356 8300 14368
rect 8352 14396 8358 14408
rect 10962 14396 10968 14408
rect 8352 14368 10968 14396
rect 8352 14356 8358 14368
rect 10962 14356 10968 14368
rect 11020 14356 11026 14408
rect 13722 14356 13728 14408
rect 13780 14396 13786 14408
rect 14277 14399 14335 14405
rect 14277 14396 14289 14399
rect 13780 14368 14289 14396
rect 13780 14356 13786 14368
rect 14277 14365 14289 14368
rect 14323 14396 14335 14399
rect 14366 14396 14372 14408
rect 14323 14368 14372 14396
rect 14323 14365 14335 14368
rect 14277 14359 14335 14365
rect 14366 14356 14372 14368
rect 14424 14356 14430 14408
rect 14476 14405 14504 14436
rect 14744 14433 14756 14467
rect 14790 14433 14802 14467
rect 14844 14464 14872 14572
rect 15013 14467 15071 14473
rect 15013 14464 15025 14467
rect 14844 14436 15025 14464
rect 14744 14427 14802 14433
rect 15013 14433 15025 14436
rect 15059 14464 15071 14467
rect 16942 14464 16948 14476
rect 15059 14436 16948 14464
rect 15059 14433 15071 14436
rect 15013 14427 15071 14433
rect 16942 14424 16948 14436
rect 17000 14424 17006 14476
rect 17310 14424 17316 14476
rect 17368 14424 17374 14476
rect 14461 14399 14519 14405
rect 14461 14365 14473 14399
rect 14507 14365 14519 14399
rect 14461 14359 14519 14365
rect 5534 14328 5540 14340
rect 4264 14300 5540 14328
rect 4157 14291 4215 14297
rect 5534 14288 5540 14300
rect 5592 14288 5598 14340
rect 14476 14328 14504 14359
rect 14642 14356 14648 14408
rect 14700 14356 14706 14408
rect 16850 14356 16856 14408
rect 16908 14396 16914 14408
rect 17037 14399 17095 14405
rect 17037 14396 17049 14399
rect 16908 14368 17049 14396
rect 16908 14356 16914 14368
rect 17037 14365 17049 14368
rect 17083 14365 17095 14399
rect 17037 14359 17095 14365
rect 14476 14300 15424 14328
rect 15396 14272 15424 14300
rect 16022 14288 16028 14340
rect 16080 14288 16086 14340
rect 18046 14288 18052 14340
rect 18104 14288 18110 14340
rect 1670 14220 1676 14272
rect 1728 14220 1734 14272
rect 1762 14220 1768 14272
rect 1820 14220 1826 14272
rect 3510 14220 3516 14272
rect 3568 14260 3574 14272
rect 4522 14260 4528 14272
rect 3568 14232 4528 14260
rect 3568 14220 3574 14232
rect 4522 14220 4528 14232
rect 4580 14220 4586 14272
rect 14185 14263 14243 14269
rect 14185 14229 14197 14263
rect 14231 14260 14243 14263
rect 14274 14260 14280 14272
rect 14231 14232 14280 14260
rect 14231 14229 14243 14232
rect 14185 14223 14243 14229
rect 14274 14220 14280 14232
rect 14332 14220 14338 14272
rect 14458 14220 14464 14272
rect 14516 14220 14522 14272
rect 15378 14220 15384 14272
rect 15436 14220 15442 14272
rect 16482 14220 16488 14272
rect 16540 14220 16546 14272
rect 18230 14220 18236 14272
rect 18288 14260 18294 14272
rect 18785 14263 18843 14269
rect 18785 14260 18797 14263
rect 18288 14232 18797 14260
rect 18288 14220 18294 14232
rect 18785 14229 18797 14232
rect 18831 14229 18843 14263
rect 18785 14223 18843 14229
rect 1104 14170 19136 14192
rect 1104 14118 3010 14170
rect 3062 14118 3074 14170
rect 3126 14118 3138 14170
rect 3190 14118 3202 14170
rect 3254 14118 3266 14170
rect 3318 14118 19136 14170
rect 1104 14096 19136 14118
rect 1670 14016 1676 14068
rect 1728 14056 1734 14068
rect 1765 14059 1823 14065
rect 1765 14056 1777 14059
rect 1728 14028 1777 14056
rect 1728 14016 1734 14028
rect 1765 14025 1777 14028
rect 1811 14025 1823 14059
rect 1765 14019 1823 14025
rect 17037 14059 17095 14065
rect 17037 14025 17049 14059
rect 17083 14056 17095 14059
rect 17402 14056 17408 14068
rect 17083 14028 17408 14056
rect 17083 14025 17095 14028
rect 17037 14019 17095 14025
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 18046 14016 18052 14068
rect 18104 14016 18110 14068
rect 18782 14016 18788 14068
rect 18840 14016 18846 14068
rect 1026 13948 1032 14000
rect 1084 13988 1090 14000
rect 1084 13960 1992 13988
rect 1084 13948 1090 13960
rect 1486 13880 1492 13932
rect 1544 13880 1550 13932
rect 1964 13929 1992 13960
rect 2682 13948 2688 14000
rect 2740 13988 2746 14000
rect 5353 13991 5411 13997
rect 2740 13960 3556 13988
rect 2740 13948 2746 13960
rect 1949 13923 2007 13929
rect 1949 13889 1961 13923
rect 1995 13889 2007 13923
rect 1949 13883 2007 13889
rect 2130 13880 2136 13932
rect 2188 13920 2194 13932
rect 3528 13929 3556 13960
rect 5353 13957 5365 13991
rect 5399 13988 5411 13991
rect 5629 13991 5687 13997
rect 5629 13988 5641 13991
rect 5399 13960 5641 13988
rect 5399 13957 5411 13960
rect 5353 13951 5411 13957
rect 5629 13957 5641 13960
rect 5675 13957 5687 13991
rect 5629 13951 5687 13957
rect 3145 13923 3203 13929
rect 3145 13920 3157 13923
rect 2188 13892 3157 13920
rect 2188 13880 2194 13892
rect 3145 13889 3157 13892
rect 3191 13889 3203 13923
rect 3145 13883 3203 13889
rect 3513 13923 3571 13929
rect 3513 13889 3525 13923
rect 3559 13889 3571 13923
rect 3513 13883 3571 13889
rect 3878 13880 3884 13932
rect 3936 13920 3942 13932
rect 4157 13923 4215 13929
rect 4157 13920 4169 13923
rect 3936 13892 4169 13920
rect 3936 13880 3942 13892
rect 4157 13889 4169 13892
rect 4203 13920 4215 13923
rect 4246 13920 4252 13932
rect 4203 13892 4252 13920
rect 4203 13889 4215 13892
rect 4157 13883 4215 13889
rect 4246 13880 4252 13892
rect 4304 13880 4310 13932
rect 4341 13923 4399 13929
rect 4341 13889 4353 13923
rect 4387 13889 4399 13923
rect 4341 13883 4399 13889
rect 3605 13855 3663 13861
rect 3605 13821 3617 13855
rect 3651 13852 3663 13855
rect 4062 13852 4068 13864
rect 3651 13824 4068 13852
rect 3651 13821 3663 13824
rect 3605 13815 3663 13821
rect 4062 13812 4068 13824
rect 4120 13852 4126 13864
rect 4356 13852 4384 13883
rect 4614 13880 4620 13932
rect 4672 13920 4678 13932
rect 4985 13923 5043 13929
rect 4985 13920 4997 13923
rect 4672 13892 4997 13920
rect 4672 13880 4678 13892
rect 4985 13889 4997 13892
rect 5031 13889 5043 13923
rect 4985 13883 5043 13889
rect 5139 13923 5197 13929
rect 5139 13889 5151 13923
rect 5185 13920 5197 13923
rect 5185 13892 5396 13920
rect 5185 13889 5197 13892
rect 5139 13883 5197 13889
rect 4120 13824 4384 13852
rect 5368 13852 5396 13892
rect 13354 13880 13360 13932
rect 13412 13880 13418 13932
rect 16574 13880 16580 13932
rect 16632 13920 16638 13932
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 16632 13892 16681 13920
rect 16632 13880 16638 13892
rect 16669 13889 16681 13892
rect 16715 13920 16727 13923
rect 16758 13920 16764 13932
rect 16715 13892 16764 13920
rect 16715 13889 16727 13892
rect 16669 13883 16727 13889
rect 16758 13880 16764 13892
rect 16816 13880 16822 13932
rect 17957 13923 18015 13929
rect 17957 13889 17969 13923
rect 18003 13920 18015 13923
rect 18414 13920 18420 13932
rect 18003 13892 18420 13920
rect 18003 13889 18015 13892
rect 17957 13883 18015 13889
rect 5368 13824 5488 13852
rect 4120 13812 4126 13824
rect 1673 13787 1731 13793
rect 1673 13753 1685 13787
rect 1719 13784 1731 13787
rect 1762 13784 1768 13796
rect 1719 13756 1768 13784
rect 1719 13753 1731 13756
rect 1673 13747 1731 13753
rect 1762 13744 1768 13756
rect 1820 13744 1826 13796
rect 5460 13784 5488 13824
rect 5534 13812 5540 13864
rect 5592 13812 5598 13864
rect 5810 13812 5816 13864
rect 5868 13812 5874 13864
rect 14366 13812 14372 13864
rect 14424 13852 14430 13864
rect 16114 13852 16120 13864
rect 14424 13824 16120 13852
rect 14424 13812 14430 13824
rect 16114 13812 16120 13824
rect 16172 13852 16178 13864
rect 17494 13852 17500 13864
rect 16172 13824 17500 13852
rect 16172 13812 16178 13824
rect 17494 13812 17500 13824
rect 17552 13852 17558 13864
rect 17972 13852 18000 13883
rect 18414 13880 18420 13892
rect 18472 13880 18478 13932
rect 18598 13880 18604 13932
rect 18656 13880 18662 13932
rect 17552 13824 18000 13852
rect 17552 13812 17558 13824
rect 5994 13784 6000 13796
rect 5460 13756 6000 13784
rect 5994 13744 6000 13756
rect 6052 13744 6058 13796
rect 3053 13719 3111 13725
rect 3053 13685 3065 13719
rect 3099 13716 3111 13719
rect 3142 13716 3148 13728
rect 3099 13688 3148 13716
rect 3099 13685 3111 13688
rect 3053 13679 3111 13685
rect 3142 13676 3148 13688
rect 3200 13676 3206 13728
rect 4341 13719 4399 13725
rect 4341 13685 4353 13719
rect 4387 13716 4399 13719
rect 4614 13716 4620 13728
rect 4387 13688 4620 13716
rect 4387 13685 4399 13688
rect 4341 13679 4399 13685
rect 4614 13676 4620 13688
rect 4672 13676 4678 13728
rect 17034 13676 17040 13728
rect 17092 13676 17098 13728
rect 17218 13676 17224 13728
rect 17276 13676 17282 13728
rect 1104 13626 19136 13648
rect 1104 13574 2350 13626
rect 2402 13574 2414 13626
rect 2466 13574 2478 13626
rect 2530 13574 2542 13626
rect 2594 13574 2606 13626
rect 2658 13574 19136 13626
rect 1104 13552 19136 13574
rect 3786 13472 3792 13524
rect 3844 13512 3850 13524
rect 5810 13512 5816 13524
rect 3844 13484 5816 13512
rect 3844 13472 3850 13484
rect 5810 13472 5816 13484
rect 5868 13472 5874 13524
rect 5994 13472 6000 13524
rect 6052 13512 6058 13524
rect 6089 13515 6147 13521
rect 6089 13512 6101 13515
rect 6052 13484 6101 13512
rect 6052 13472 6058 13484
rect 6089 13481 6101 13484
rect 6135 13481 6147 13515
rect 6089 13475 6147 13481
rect 13906 13472 13912 13524
rect 13964 13512 13970 13524
rect 15102 13512 15108 13524
rect 13964 13484 15108 13512
rect 13964 13472 13970 13484
rect 15102 13472 15108 13484
rect 15160 13512 15166 13524
rect 15381 13515 15439 13521
rect 15381 13512 15393 13515
rect 15160 13484 15393 13512
rect 15160 13472 15166 13484
rect 15381 13481 15393 13484
rect 15427 13481 15439 13515
rect 15381 13475 15439 13481
rect 16022 13472 16028 13524
rect 16080 13472 16086 13524
rect 18598 13472 18604 13524
rect 18656 13472 18662 13524
rect 13648 13416 15884 13444
rect 1854 13336 1860 13388
rect 1912 13376 1918 13388
rect 4341 13379 4399 13385
rect 4341 13376 4353 13379
rect 1912 13348 4353 13376
rect 1912 13336 1918 13348
rect 4341 13345 4353 13348
rect 4387 13345 4399 13379
rect 4341 13339 4399 13345
rect 4614 13336 4620 13388
rect 4672 13336 4678 13388
rect 1765 13311 1823 13317
rect 1765 13277 1777 13311
rect 1811 13308 1823 13311
rect 1811 13280 1900 13308
rect 1811 13277 1823 13280
rect 1765 13271 1823 13277
rect 1578 13132 1584 13184
rect 1636 13132 1642 13184
rect 1872 13172 1900 13280
rect 4062 13268 4068 13320
rect 4120 13268 4126 13320
rect 4249 13311 4307 13317
rect 4249 13277 4261 13311
rect 4295 13277 4307 13311
rect 4249 13271 4307 13277
rect 2130 13200 2136 13252
rect 2188 13200 2194 13252
rect 3142 13200 3148 13252
rect 3200 13200 3206 13252
rect 3878 13200 3884 13252
rect 3936 13240 3942 13252
rect 4264 13240 4292 13271
rect 6362 13268 6368 13320
rect 6420 13308 6426 13320
rect 6638 13308 6644 13320
rect 6420 13280 6644 13308
rect 6420 13268 6426 13280
rect 6638 13268 6644 13280
rect 6696 13268 6702 13320
rect 13648 13317 13676 13416
rect 14458 13376 14464 13388
rect 13832 13348 14464 13376
rect 13832 13317 13860 13348
rect 14458 13336 14464 13348
rect 14516 13336 14522 13388
rect 15856 13376 15884 13416
rect 16577 13379 16635 13385
rect 16577 13376 16589 13379
rect 15856 13348 16589 13376
rect 16577 13345 16589 13348
rect 16623 13376 16635 13379
rect 17218 13376 17224 13388
rect 16623 13348 17224 13376
rect 16623 13345 16635 13348
rect 16577 13339 16635 13345
rect 17218 13336 17224 13348
rect 17276 13336 17282 13388
rect 18049 13379 18107 13385
rect 18049 13345 18061 13379
rect 18095 13376 18107 13379
rect 18095 13348 18460 13376
rect 18095 13345 18107 13348
rect 18049 13339 18107 13345
rect 13633 13311 13691 13317
rect 13633 13277 13645 13311
rect 13679 13277 13691 13311
rect 13633 13271 13691 13277
rect 13817 13311 13875 13317
rect 13817 13277 13829 13311
rect 13863 13277 13875 13311
rect 13817 13271 13875 13277
rect 13909 13311 13967 13317
rect 13909 13277 13921 13311
rect 13955 13308 13967 13311
rect 13998 13308 14004 13320
rect 13955 13280 14004 13308
rect 13955 13277 13967 13280
rect 13909 13271 13967 13277
rect 13998 13268 14004 13280
rect 14056 13268 14062 13320
rect 14093 13311 14151 13317
rect 14093 13277 14105 13311
rect 14139 13308 14151 13311
rect 14182 13308 14188 13320
rect 14139 13280 14188 13308
rect 14139 13277 14151 13280
rect 14093 13271 14151 13277
rect 6273 13243 6331 13249
rect 6273 13240 6285 13243
rect 3936 13212 4292 13240
rect 5842 13212 6285 13240
rect 3936 13200 3942 13212
rect 6273 13209 6285 13212
rect 6319 13209 6331 13243
rect 6273 13203 6331 13209
rect 10962 13200 10968 13252
rect 11020 13240 11026 13252
rect 14108 13240 14136 13271
rect 14182 13268 14188 13280
rect 14240 13268 14246 13320
rect 15746 13268 15752 13320
rect 15804 13308 15810 13320
rect 16114 13308 16120 13320
rect 15804 13280 16120 13308
rect 15804 13268 15810 13280
rect 16114 13268 16120 13280
rect 16172 13268 16178 13320
rect 18432 13317 18460 13348
rect 16301 13311 16359 13317
rect 16301 13277 16313 13311
rect 16347 13277 16359 13311
rect 16301 13271 16359 13277
rect 18325 13311 18383 13317
rect 18325 13277 18337 13311
rect 18371 13277 18383 13311
rect 18325 13271 18383 13277
rect 18417 13311 18475 13317
rect 18417 13277 18429 13311
rect 18463 13277 18475 13311
rect 18417 13271 18475 13277
rect 11020 13212 14136 13240
rect 11020 13200 11026 13212
rect 15102 13200 15108 13252
rect 15160 13240 15166 13252
rect 16316 13240 16344 13271
rect 16850 13240 16856 13252
rect 15160 13212 16856 13240
rect 15160 13200 15166 13212
rect 16850 13200 16856 13212
rect 16908 13200 16914 13252
rect 18233 13243 18291 13249
rect 18233 13240 18245 13243
rect 17802 13212 18245 13240
rect 18233 13209 18245 13212
rect 18279 13209 18291 13243
rect 18340 13240 18368 13271
rect 18340 13212 18460 13240
rect 18233 13203 18291 13209
rect 18432 13184 18460 13212
rect 2866 13172 2872 13184
rect 1872 13144 2872 13172
rect 2866 13132 2872 13144
rect 2924 13172 2930 13184
rect 3605 13175 3663 13181
rect 3605 13172 3617 13175
rect 2924 13144 3617 13172
rect 2924 13132 2930 13144
rect 3605 13141 3617 13144
rect 3651 13141 3663 13175
rect 3605 13135 3663 13141
rect 3970 13132 3976 13184
rect 4028 13132 4034 13184
rect 13170 13132 13176 13184
rect 13228 13172 13234 13184
rect 13449 13175 13507 13181
rect 13449 13172 13461 13175
rect 13228 13144 13461 13172
rect 13228 13132 13234 13144
rect 13449 13141 13461 13144
rect 13495 13141 13507 13175
rect 13449 13135 13507 13141
rect 18414 13132 18420 13184
rect 18472 13132 18478 13184
rect 1104 13082 19136 13104
rect 1104 13030 3010 13082
rect 3062 13030 3074 13082
rect 3126 13030 3138 13082
rect 3190 13030 3202 13082
rect 3254 13030 3266 13082
rect 3318 13030 19136 13082
rect 1104 13008 19136 13030
rect 1210 12928 1216 12980
rect 1268 12968 1274 12980
rect 1397 12971 1455 12977
rect 1397 12968 1409 12971
rect 1268 12940 1409 12968
rect 1268 12928 1274 12940
rect 1397 12937 1409 12940
rect 1443 12937 1455 12971
rect 1397 12931 1455 12937
rect 2130 12928 2136 12980
rect 2188 12968 2194 12980
rect 2593 12971 2651 12977
rect 2593 12968 2605 12971
rect 2188 12940 2605 12968
rect 2188 12928 2194 12940
rect 2593 12937 2605 12940
rect 2639 12937 2651 12971
rect 2593 12931 2651 12937
rect 13354 12928 13360 12980
rect 13412 12968 13418 12980
rect 13906 12968 13912 12980
rect 13412 12940 13912 12968
rect 13412 12928 13418 12940
rect 13906 12928 13912 12940
rect 13964 12928 13970 12980
rect 13998 12928 14004 12980
rect 14056 12968 14062 12980
rect 14645 12971 14703 12977
rect 14645 12968 14657 12971
rect 14056 12940 14657 12968
rect 14056 12928 14062 12940
rect 14645 12937 14657 12940
rect 14691 12968 14703 12971
rect 15470 12968 15476 12980
rect 14691 12940 15476 12968
rect 14691 12937 14703 12940
rect 14645 12931 14703 12937
rect 15470 12928 15476 12940
rect 15528 12928 15534 12980
rect 15654 12928 15660 12980
rect 15712 12928 15718 12980
rect 18322 12928 18328 12980
rect 18380 12928 18386 12980
rect 18506 12928 18512 12980
rect 18564 12968 18570 12980
rect 18601 12971 18659 12977
rect 18601 12968 18613 12971
rect 18564 12940 18613 12968
rect 18564 12928 18570 12940
rect 18601 12937 18613 12940
rect 18647 12937 18659 12971
rect 18601 12931 18659 12937
rect 3418 12900 3424 12912
rect 3068 12872 3424 12900
rect 1578 12792 1584 12844
rect 1636 12792 1642 12844
rect 1670 12792 1676 12844
rect 1728 12792 1734 12844
rect 1762 12792 1768 12844
rect 1820 12832 1826 12844
rect 2777 12835 2835 12841
rect 2777 12832 2789 12835
rect 1820 12804 2789 12832
rect 1820 12792 1826 12804
rect 2777 12801 2789 12804
rect 2823 12801 2835 12835
rect 2777 12795 2835 12801
rect 2866 12792 2872 12844
rect 2924 12792 2930 12844
rect 3068 12841 3096 12872
rect 3418 12860 3424 12872
rect 3476 12900 3482 12912
rect 5350 12900 5356 12912
rect 3476 12872 5356 12900
rect 3476 12860 3482 12872
rect 5350 12860 5356 12872
rect 5408 12860 5414 12912
rect 13372 12900 13400 12928
rect 12912 12872 13400 12900
rect 3053 12835 3111 12841
rect 3053 12801 3065 12835
rect 3099 12801 3111 12835
rect 3053 12795 3111 12801
rect 3237 12835 3295 12841
rect 3237 12801 3249 12835
rect 3283 12832 3295 12835
rect 3970 12832 3976 12844
rect 3283 12804 3976 12832
rect 3283 12801 3295 12804
rect 3237 12795 3295 12801
rect 3970 12792 3976 12804
rect 4028 12792 4034 12844
rect 12912 12841 12940 12872
rect 12897 12835 12955 12841
rect 12897 12801 12909 12835
rect 12943 12801 12955 12835
rect 12897 12795 12955 12801
rect 14274 12792 14280 12844
rect 14332 12792 14338 12844
rect 15194 12792 15200 12844
rect 15252 12832 15258 12844
rect 15289 12835 15347 12841
rect 15289 12832 15301 12835
rect 15252 12804 15301 12832
rect 15252 12792 15258 12804
rect 15289 12801 15301 12804
rect 15335 12801 15347 12835
rect 15289 12795 15347 12801
rect 15443 12835 15501 12841
rect 15443 12801 15455 12835
rect 15489 12832 15501 12835
rect 16482 12832 16488 12844
rect 15489 12804 16488 12832
rect 15489 12801 15501 12804
rect 15443 12795 15501 12801
rect 16482 12792 16488 12804
rect 16540 12792 16546 12844
rect 18138 12792 18144 12844
rect 18196 12792 18202 12844
rect 18782 12792 18788 12844
rect 18840 12792 18846 12844
rect 2961 12767 3019 12773
rect 2961 12733 2973 12767
rect 3007 12764 3019 12767
rect 4062 12764 4068 12776
rect 3007 12736 4068 12764
rect 3007 12733 3019 12736
rect 2961 12727 3019 12733
rect 4062 12724 4068 12736
rect 4120 12724 4126 12776
rect 13170 12724 13176 12776
rect 13228 12724 13234 12776
rect 1857 12631 1915 12637
rect 1857 12597 1869 12631
rect 1903 12628 1915 12631
rect 7006 12628 7012 12640
rect 1903 12600 7012 12628
rect 1903 12597 1915 12600
rect 1857 12591 1915 12597
rect 7006 12588 7012 12600
rect 7064 12588 7070 12640
rect 1104 12538 19136 12560
rect 1104 12486 2350 12538
rect 2402 12486 2414 12538
rect 2466 12486 2478 12538
rect 2530 12486 2542 12538
rect 2594 12486 2606 12538
rect 2658 12486 19136 12538
rect 1104 12464 19136 12486
rect 11882 12384 11888 12436
rect 11940 12424 11946 12436
rect 15102 12424 15108 12436
rect 11940 12396 15108 12424
rect 11940 12384 11946 12396
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 13906 12248 13912 12300
rect 13964 12288 13970 12300
rect 14093 12291 14151 12297
rect 14093 12288 14105 12291
rect 13964 12260 14105 12288
rect 13964 12248 13970 12260
rect 14093 12257 14105 12260
rect 14139 12257 14151 12291
rect 14093 12251 14151 12257
rect 18048 12223 18106 12229
rect 18048 12189 18060 12223
rect 18094 12189 18106 12223
rect 18048 12183 18106 12189
rect 11882 12112 11888 12164
rect 11940 12112 11946 12164
rect 12986 12112 12992 12164
rect 13044 12112 13050 12164
rect 13633 12155 13691 12161
rect 13633 12121 13645 12155
rect 13679 12121 13691 12155
rect 13633 12115 13691 12121
rect 3878 12044 3884 12096
rect 3936 12084 3942 12096
rect 4430 12084 4436 12096
rect 3936 12056 4436 12084
rect 3936 12044 3942 12056
rect 4430 12044 4436 12056
rect 4488 12044 4494 12096
rect 13648 12084 13676 12115
rect 14366 12112 14372 12164
rect 14424 12112 14430 12164
rect 15102 12112 15108 12164
rect 15160 12112 15166 12164
rect 17402 12112 17408 12164
rect 17460 12152 17466 12164
rect 18064 12152 18092 12183
rect 18138 12180 18144 12232
rect 18196 12220 18202 12232
rect 18690 12220 18696 12232
rect 18196 12192 18696 12220
rect 18196 12180 18202 12192
rect 18690 12180 18696 12192
rect 18748 12180 18754 12232
rect 18782 12180 18788 12232
rect 18840 12180 18846 12232
rect 17460 12124 18644 12152
rect 17460 12112 17466 12124
rect 15378 12084 15384 12096
rect 13648 12056 15384 12084
rect 15378 12044 15384 12056
rect 15436 12044 15442 12096
rect 15654 12044 15660 12096
rect 15712 12084 15718 12096
rect 15841 12087 15899 12093
rect 15841 12084 15853 12087
rect 15712 12056 15853 12084
rect 15712 12044 15718 12056
rect 15841 12053 15853 12056
rect 15887 12053 15899 12087
rect 15841 12047 15899 12053
rect 17586 12044 17592 12096
rect 17644 12084 17650 12096
rect 18616 12093 18644 12124
rect 17773 12087 17831 12093
rect 17773 12084 17785 12087
rect 17644 12056 17785 12084
rect 17644 12044 17650 12056
rect 17773 12053 17785 12056
rect 17819 12053 17831 12087
rect 17773 12047 17831 12053
rect 18601 12087 18659 12093
rect 18601 12053 18613 12087
rect 18647 12053 18659 12087
rect 18601 12047 18659 12053
rect 1104 11994 19136 12016
rect 1104 11942 3010 11994
rect 3062 11942 3074 11994
rect 3126 11942 3138 11994
rect 3190 11942 3202 11994
rect 3254 11942 3266 11994
rect 3318 11942 19136 11994
rect 1104 11920 19136 11942
rect 1780 11852 3280 11880
rect 1780 11824 1808 11852
rect 1673 11815 1731 11821
rect 1673 11781 1685 11815
rect 1719 11812 1731 11815
rect 1762 11812 1768 11824
rect 1719 11784 1768 11812
rect 1719 11781 1731 11784
rect 1673 11775 1731 11781
rect 1762 11772 1768 11784
rect 1820 11772 1826 11824
rect 2130 11772 2136 11824
rect 2188 11772 2194 11824
rect 3252 11744 3280 11852
rect 4154 11840 4160 11892
rect 4212 11880 4218 11892
rect 4798 11880 4804 11892
rect 4212 11852 4804 11880
rect 4212 11840 4218 11852
rect 4798 11840 4804 11852
rect 4856 11840 4862 11892
rect 12986 11840 12992 11892
rect 13044 11840 13050 11892
rect 15102 11840 15108 11892
rect 15160 11840 15166 11892
rect 18690 11840 18696 11892
rect 18748 11840 18754 11892
rect 4356 11784 5028 11812
rect 3878 11744 3884 11756
rect 3252 11716 3884 11744
rect 3878 11704 3884 11716
rect 3936 11744 3942 11756
rect 3973 11747 4031 11753
rect 3973 11744 3985 11747
rect 3936 11716 3985 11744
rect 3936 11704 3942 11716
rect 3973 11713 3985 11716
rect 4019 11713 4031 11747
rect 3973 11707 4031 11713
rect 4062 11704 4068 11756
rect 4120 11704 4126 11756
rect 4154 11704 4160 11756
rect 4212 11704 4218 11756
rect 4356 11753 4384 11784
rect 5000 11756 5028 11784
rect 5074 11772 5080 11824
rect 5132 11812 5138 11824
rect 9309 11815 9367 11821
rect 9309 11812 9321 11815
rect 5132 11784 9321 11812
rect 5132 11772 5138 11784
rect 9309 11781 9321 11784
rect 9355 11781 9367 11815
rect 9309 11775 9367 11781
rect 16485 11815 16543 11821
rect 16485 11781 16497 11815
rect 16531 11812 16543 11815
rect 17494 11812 17500 11824
rect 16531 11784 17500 11812
rect 16531 11781 16543 11784
rect 16485 11775 16543 11781
rect 17494 11772 17500 11784
rect 17552 11772 17558 11824
rect 17954 11772 17960 11824
rect 18012 11772 18018 11824
rect 4341 11747 4399 11753
rect 4341 11713 4353 11747
rect 4387 11713 4399 11747
rect 4341 11707 4399 11713
rect 4430 11704 4436 11756
rect 4488 11704 4494 11756
rect 4798 11704 4804 11756
rect 4856 11704 4862 11756
rect 4982 11704 4988 11756
rect 5040 11704 5046 11756
rect 5445 11747 5503 11753
rect 5445 11713 5457 11747
rect 5491 11744 5503 11747
rect 6362 11744 6368 11756
rect 5491 11716 6368 11744
rect 5491 11713 5503 11716
rect 5445 11707 5503 11713
rect 6362 11704 6368 11716
rect 6420 11704 6426 11756
rect 13081 11747 13139 11753
rect 13081 11713 13093 11747
rect 13127 11744 13139 11747
rect 15013 11747 15071 11753
rect 15013 11744 15025 11747
rect 13127 11716 15025 11744
rect 13127 11713 13139 11716
rect 13081 11707 13139 11713
rect 15013 11713 15025 11716
rect 15059 11744 15071 11747
rect 15059 11716 15148 11744
rect 15059 11713 15071 11716
rect 15013 11707 15071 11713
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 1762 11676 1768 11688
rect 1443 11648 1768 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 1762 11636 1768 11648
rect 1820 11636 1826 11688
rect 4080 11676 4108 11704
rect 4080 11648 4292 11676
rect 3142 11500 3148 11552
rect 3200 11500 3206 11552
rect 3697 11543 3755 11549
rect 3697 11509 3709 11543
rect 3743 11540 3755 11543
rect 4154 11540 4160 11552
rect 3743 11512 4160 11540
rect 3743 11509 3755 11512
rect 3697 11503 3755 11509
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 4264 11540 4292 11648
rect 4706 11636 4712 11688
rect 4764 11636 4770 11688
rect 4525 11543 4583 11549
rect 4525 11540 4537 11543
rect 4264 11512 4537 11540
rect 4525 11509 4537 11512
rect 4571 11509 4583 11543
rect 4525 11503 4583 11509
rect 4890 11500 4896 11552
rect 4948 11500 4954 11552
rect 5074 11500 5080 11552
rect 5132 11500 5138 11552
rect 5258 11500 5264 11552
rect 5316 11540 5322 11552
rect 5353 11543 5411 11549
rect 5353 11540 5365 11543
rect 5316 11512 5365 11540
rect 5316 11500 5322 11512
rect 5353 11509 5365 11512
rect 5399 11509 5411 11543
rect 5353 11503 5411 11509
rect 10594 11500 10600 11552
rect 10652 11540 10658 11552
rect 10962 11540 10968 11552
rect 10652 11512 10968 11540
rect 10652 11500 10658 11512
rect 10962 11500 10968 11512
rect 11020 11500 11026 11552
rect 15120 11540 15148 11716
rect 15194 11704 15200 11756
rect 15252 11744 15258 11756
rect 15381 11747 15439 11753
rect 15381 11744 15393 11747
rect 15252 11716 15393 11744
rect 15252 11704 15258 11716
rect 15381 11713 15393 11716
rect 15427 11713 15439 11747
rect 15381 11707 15439 11713
rect 15535 11747 15593 11753
rect 15535 11713 15547 11747
rect 15581 11744 15593 11747
rect 15654 11744 15660 11756
rect 15581 11716 15660 11744
rect 15581 11713 15593 11716
rect 15535 11707 15593 11713
rect 15396 11608 15424 11707
rect 15654 11704 15660 11716
rect 15712 11704 15718 11756
rect 15749 11747 15807 11753
rect 15749 11713 15761 11747
rect 15795 11744 15807 11747
rect 16025 11747 16083 11753
rect 16025 11744 16037 11747
rect 15795 11716 16037 11744
rect 15795 11713 15807 11716
rect 15749 11707 15807 11713
rect 16025 11713 16037 11716
rect 16071 11713 16083 11747
rect 16025 11707 16083 11713
rect 16942 11704 16948 11756
rect 17000 11704 17006 11756
rect 15838 11636 15844 11688
rect 15896 11636 15902 11688
rect 17218 11636 17224 11688
rect 17276 11636 17282 11688
rect 15930 11608 15936 11620
rect 15396 11580 15936 11608
rect 15930 11568 15936 11580
rect 15988 11568 15994 11620
rect 15746 11540 15752 11552
rect 15120 11512 15752 11540
rect 15746 11500 15752 11512
rect 15804 11500 15810 11552
rect 1104 11450 19136 11472
rect 1104 11398 2350 11450
rect 2402 11398 2414 11450
rect 2466 11398 2478 11450
rect 2530 11398 2542 11450
rect 2594 11398 2606 11450
rect 2658 11398 19136 11450
rect 1104 11376 19136 11398
rect 2130 11296 2136 11348
rect 2188 11296 2194 11348
rect 3237 11339 3295 11345
rect 3237 11305 3249 11339
rect 3283 11336 3295 11339
rect 4062 11336 4068 11348
rect 3283 11308 4068 11336
rect 3283 11305 3295 11308
rect 3237 11299 3295 11305
rect 4062 11296 4068 11308
rect 4120 11296 4126 11348
rect 4341 11339 4399 11345
rect 4341 11305 4353 11339
rect 4387 11336 4399 11339
rect 4706 11336 4712 11348
rect 4387 11308 4712 11336
rect 4387 11305 4399 11308
rect 4341 11299 4399 11305
rect 4706 11296 4712 11308
rect 4764 11296 4770 11348
rect 5169 11339 5227 11345
rect 5169 11305 5181 11339
rect 5215 11305 5227 11339
rect 5169 11299 5227 11305
rect 5261 11339 5319 11345
rect 5261 11305 5273 11339
rect 5307 11336 5319 11339
rect 5350 11336 5356 11348
rect 5307 11308 5356 11336
rect 5307 11305 5319 11308
rect 5261 11299 5319 11305
rect 3142 11228 3148 11280
rect 3200 11228 3206 11280
rect 3786 11228 3792 11280
rect 3844 11268 3850 11280
rect 4798 11268 4804 11280
rect 3844 11240 4804 11268
rect 3844 11228 3850 11240
rect 3513 11203 3571 11209
rect 3513 11169 3525 11203
rect 3559 11200 3571 11203
rect 3559 11172 4108 11200
rect 3559 11169 3571 11172
rect 3513 11163 3571 11169
rect 1394 11092 1400 11144
rect 1452 11092 1458 11144
rect 2222 11092 2228 11144
rect 2280 11092 2286 11144
rect 3605 11135 3663 11141
rect 3605 11101 3617 11135
rect 3651 11132 3663 11135
rect 3651 11104 3832 11132
rect 3651 11101 3663 11104
rect 3605 11095 3663 11101
rect 2774 11024 2780 11076
rect 2832 11064 2838 11076
rect 3510 11064 3516 11076
rect 2832 11036 3516 11064
rect 2832 11024 2838 11036
rect 3510 11024 3516 11036
rect 3568 11024 3574 11076
rect 1578 10956 1584 11008
rect 1636 10956 1642 11008
rect 3804 10996 3832 11104
rect 3878 11092 3884 11144
rect 3936 11092 3942 11144
rect 4080 11064 4108 11172
rect 4172 11141 4200 11240
rect 4798 11228 4804 11240
rect 4856 11228 4862 11280
rect 4890 11228 4896 11280
rect 4948 11268 4954 11280
rect 5184 11268 5212 11299
rect 5350 11296 5356 11308
rect 5408 11296 5414 11348
rect 5534 11296 5540 11348
rect 5592 11296 5598 11348
rect 6362 11296 6368 11348
rect 6420 11336 6426 11348
rect 16577 11339 16635 11345
rect 16577 11336 16589 11339
rect 6420 11308 7604 11336
rect 6420 11296 6426 11308
rect 5552 11268 5580 11296
rect 4948 11240 5120 11268
rect 5184 11240 5580 11268
rect 4948 11228 4954 11240
rect 4709 11203 4767 11209
rect 4709 11169 4721 11203
rect 4755 11200 4767 11203
rect 4985 11203 5043 11209
rect 4985 11200 4997 11203
rect 4755 11172 4997 11200
rect 4755 11169 4767 11172
rect 4709 11163 4767 11169
rect 4985 11169 4997 11172
rect 5031 11169 5043 11203
rect 5092 11200 5120 11240
rect 5169 11203 5227 11209
rect 5169 11200 5181 11203
rect 5092 11172 5181 11200
rect 4985 11163 5043 11169
rect 5169 11169 5181 11172
rect 5215 11169 5227 11203
rect 5169 11163 5227 11169
rect 5537 11203 5595 11209
rect 5537 11169 5549 11203
rect 5583 11200 5595 11203
rect 5810 11200 5816 11212
rect 5583 11172 5816 11200
rect 5583 11169 5595 11172
rect 5537 11163 5595 11169
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 6822 11160 6828 11212
rect 6880 11200 6886 11212
rect 7285 11203 7343 11209
rect 7285 11200 7297 11203
rect 6880 11172 7297 11200
rect 6880 11160 6886 11172
rect 7285 11169 7297 11172
rect 7331 11169 7343 11203
rect 7285 11163 7343 11169
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11101 4215 11135
rect 4157 11095 4215 11101
rect 4246 11092 4252 11144
rect 4304 11132 4310 11144
rect 4433 11135 4491 11141
rect 4433 11132 4445 11135
rect 4304 11104 4445 11132
rect 4304 11092 4310 11104
rect 4433 11101 4445 11104
rect 4479 11101 4491 11135
rect 4433 11095 4491 11101
rect 4890 11092 4896 11144
rect 4948 11092 4954 11144
rect 5074 11092 5080 11144
rect 5132 11132 5138 11144
rect 7576 11141 7604 11308
rect 15304 11308 16589 11336
rect 5353 11135 5411 11141
rect 5353 11132 5365 11135
rect 5132 11104 5365 11132
rect 5132 11092 5138 11104
rect 5353 11101 5365 11104
rect 5399 11101 5411 11135
rect 5353 11095 5411 11101
rect 7561 11135 7619 11141
rect 7561 11101 7573 11135
rect 7607 11101 7619 11135
rect 7561 11095 7619 11101
rect 14366 11092 14372 11144
rect 14424 11132 14430 11144
rect 15304 11141 15332 11308
rect 16577 11305 16589 11308
rect 16623 11305 16635 11339
rect 16577 11299 16635 11305
rect 17129 11339 17187 11345
rect 17129 11305 17141 11339
rect 17175 11336 17187 11339
rect 17218 11336 17224 11348
rect 17175 11308 17224 11336
rect 17175 11305 17187 11308
rect 17129 11299 17187 11305
rect 15378 11228 15384 11280
rect 15436 11268 15442 11280
rect 16209 11271 16267 11277
rect 16209 11268 16221 11271
rect 15436 11240 16221 11268
rect 15436 11228 15442 11240
rect 16209 11237 16221 11240
rect 16255 11268 16267 11271
rect 16482 11268 16488 11280
rect 16255 11240 16488 11268
rect 16255 11237 16267 11240
rect 16209 11231 16267 11237
rect 16482 11228 16488 11240
rect 16540 11228 16546 11280
rect 16592 11268 16620 11299
rect 17218 11296 17224 11308
rect 17276 11296 17282 11348
rect 17954 11296 17960 11348
rect 18012 11336 18018 11348
rect 18049 11339 18107 11345
rect 18049 11336 18061 11339
rect 18012 11308 18061 11336
rect 18012 11296 18018 11308
rect 18049 11305 18061 11308
rect 18095 11305 18107 11339
rect 18049 11299 18107 11305
rect 17402 11268 17408 11280
rect 16592 11240 17408 11268
rect 17402 11228 17408 11240
rect 17460 11228 17466 11280
rect 15580 11172 17816 11200
rect 15580 11144 15608 11172
rect 17788 11144 17816 11172
rect 15289 11135 15347 11141
rect 15289 11132 15301 11135
rect 14424 11104 15301 11132
rect 14424 11092 14430 11104
rect 15289 11101 15301 11104
rect 15335 11101 15347 11135
rect 15289 11095 15347 11101
rect 15473 11135 15531 11141
rect 15473 11101 15485 11135
rect 15519 11132 15531 11135
rect 15562 11132 15568 11144
rect 15519 11104 15568 11132
rect 15519 11101 15531 11104
rect 15473 11095 15531 11101
rect 15562 11092 15568 11104
rect 15620 11092 15626 11144
rect 15746 11092 15752 11144
rect 15804 11092 15810 11144
rect 17402 11092 17408 11144
rect 17460 11092 17466 11144
rect 17494 11092 17500 11144
rect 17552 11092 17558 11144
rect 17586 11092 17592 11144
rect 17644 11092 17650 11144
rect 17770 11092 17776 11144
rect 17828 11092 17834 11144
rect 17957 11135 18015 11141
rect 17957 11101 17969 11135
rect 18003 11132 18015 11135
rect 18414 11132 18420 11144
rect 18003 11104 18420 11132
rect 18003 11101 18015 11104
rect 17957 11095 18015 11101
rect 18414 11092 18420 11104
rect 18472 11092 18478 11144
rect 18782 11092 18788 11144
rect 18840 11092 18846 11144
rect 4525 11067 4583 11073
rect 4525 11064 4537 11067
rect 4080 11036 4537 11064
rect 4525 11033 4537 11036
rect 4571 11033 4583 11067
rect 5813 11067 5871 11073
rect 4525 11027 4583 11033
rect 4632 11036 5580 11064
rect 3973 10999 4031 11005
rect 3973 10996 3985 10999
rect 3804 10968 3985 10996
rect 3973 10965 3985 10968
rect 4019 10996 4031 10999
rect 4632 10996 4660 11036
rect 4019 10968 4660 10996
rect 5552 10996 5580 11036
rect 5813 11033 5825 11067
rect 5859 11064 5871 11067
rect 6086 11064 6092 11076
rect 5859 11036 6092 11064
rect 5859 11033 5871 11036
rect 5813 11027 5871 11033
rect 6086 11024 6092 11036
rect 6144 11024 6150 11076
rect 7469 11067 7527 11073
rect 7469 11064 7481 11067
rect 7038 11036 7481 11064
rect 7469 11033 7481 11036
rect 7515 11033 7527 11067
rect 7469 11027 7527 11033
rect 15654 11024 15660 11076
rect 15712 11024 15718 11076
rect 16577 11067 16635 11073
rect 16577 11033 16589 11067
rect 16623 11064 16635 11067
rect 16623 11036 18644 11064
rect 16623 11033 16635 11036
rect 16577 11027 16635 11033
rect 6822 10996 6828 11008
rect 5552 10968 6828 10996
rect 4019 10965 4031 10968
rect 3973 10959 4031 10965
rect 6822 10956 6828 10968
rect 6880 10956 6886 11008
rect 15470 10956 15476 11008
rect 15528 10956 15534 11008
rect 16761 10999 16819 11005
rect 16761 10965 16773 10999
rect 16807 10996 16819 10999
rect 16850 10996 16856 11008
rect 16807 10968 16856 10996
rect 16807 10965 16819 10968
rect 16761 10959 16819 10965
rect 16850 10956 16856 10968
rect 16908 10956 16914 11008
rect 18616 11005 18644 11036
rect 18601 10999 18659 11005
rect 18601 10965 18613 10999
rect 18647 10965 18659 10999
rect 18601 10959 18659 10965
rect 1104 10906 19136 10928
rect 1104 10854 3010 10906
rect 3062 10854 3074 10906
rect 3126 10854 3138 10906
rect 3190 10854 3202 10906
rect 3254 10854 3266 10906
rect 3318 10854 19136 10906
rect 1104 10832 19136 10854
rect 3145 10795 3203 10801
rect 3145 10761 3157 10795
rect 3191 10792 3203 10795
rect 3878 10792 3884 10804
rect 3191 10764 3884 10792
rect 3191 10761 3203 10764
rect 3145 10755 3203 10761
rect 3878 10752 3884 10764
rect 3936 10792 3942 10804
rect 4522 10792 4528 10804
rect 3936 10764 4528 10792
rect 3936 10752 3942 10764
rect 4522 10752 4528 10764
rect 4580 10752 4586 10804
rect 4890 10752 4896 10804
rect 4948 10792 4954 10804
rect 4948 10764 5672 10792
rect 4948 10752 4954 10764
rect 1578 10684 1584 10736
rect 1636 10724 1642 10736
rect 1673 10727 1731 10733
rect 1673 10724 1685 10727
rect 1636 10696 1685 10724
rect 1636 10684 1642 10696
rect 1673 10693 1685 10696
rect 1719 10693 1731 10727
rect 1673 10687 1731 10693
rect 2222 10684 2228 10736
rect 2280 10684 2286 10736
rect 5258 10724 5264 10736
rect 5106 10696 5264 10724
rect 5258 10684 5264 10696
rect 5316 10684 5322 10736
rect 5534 10684 5540 10736
rect 5592 10684 5598 10736
rect 5644 10724 5672 10764
rect 6086 10752 6092 10804
rect 6144 10792 6150 10804
rect 6365 10795 6423 10801
rect 6365 10792 6377 10795
rect 6144 10764 6377 10792
rect 6144 10752 6150 10764
rect 6365 10761 6377 10764
rect 6411 10761 6423 10795
rect 6365 10755 6423 10761
rect 6822 10752 6828 10804
rect 6880 10752 6886 10804
rect 15838 10752 15844 10804
rect 15896 10792 15902 10804
rect 16025 10795 16083 10801
rect 16025 10792 16037 10795
rect 15896 10764 16037 10792
rect 15896 10752 15902 10764
rect 16025 10761 16037 10764
rect 16071 10761 16083 10795
rect 16025 10755 16083 10761
rect 6733 10727 6791 10733
rect 6733 10724 6745 10727
rect 5644 10696 6745 10724
rect 6733 10693 6745 10696
rect 6779 10693 6791 10727
rect 6733 10687 6791 10693
rect 5810 10616 5816 10668
rect 5868 10616 5874 10668
rect 15654 10616 15660 10668
rect 15712 10616 15718 10668
rect 18141 10659 18199 10665
rect 18141 10625 18153 10659
rect 18187 10656 18199 10659
rect 18322 10656 18328 10668
rect 18187 10628 18328 10656
rect 18187 10625 18199 10628
rect 18141 10619 18199 10625
rect 18322 10616 18328 10628
rect 18380 10616 18386 10668
rect 18601 10659 18659 10665
rect 18601 10625 18613 10659
rect 18647 10625 18659 10659
rect 18601 10619 18659 10625
rect 1394 10548 1400 10600
rect 1452 10548 1458 10600
rect 4065 10591 4123 10597
rect 4065 10557 4077 10591
rect 4111 10588 4123 10591
rect 4982 10588 4988 10600
rect 4111 10560 4988 10588
rect 4111 10557 4123 10560
rect 4065 10551 4123 10557
rect 4982 10548 4988 10560
rect 5040 10548 5046 10600
rect 6730 10548 6736 10600
rect 6788 10588 6794 10600
rect 6917 10591 6975 10597
rect 6917 10588 6929 10591
rect 6788 10560 6929 10588
rect 6788 10548 6794 10560
rect 6917 10557 6929 10560
rect 6963 10557 6975 10591
rect 6917 10551 6975 10557
rect 14182 10548 14188 10600
rect 14240 10588 14246 10600
rect 14277 10591 14335 10597
rect 14277 10588 14289 10591
rect 14240 10560 14289 10588
rect 14240 10548 14246 10560
rect 14277 10557 14289 10560
rect 14323 10557 14335 10591
rect 14277 10551 14335 10557
rect 14553 10591 14611 10597
rect 14553 10557 14565 10591
rect 14599 10588 14611 10591
rect 15194 10588 15200 10600
rect 14599 10560 15200 10588
rect 14599 10557 14611 10560
rect 14553 10551 14611 10557
rect 15194 10548 15200 10560
rect 15252 10548 15258 10600
rect 17954 10548 17960 10600
rect 18012 10588 18018 10600
rect 18616 10588 18644 10619
rect 18012 10560 18644 10588
rect 18012 10548 18018 10560
rect 18325 10455 18383 10461
rect 18325 10421 18337 10455
rect 18371 10452 18383 10455
rect 18598 10452 18604 10464
rect 18371 10424 18604 10452
rect 18371 10421 18383 10424
rect 18325 10415 18383 10421
rect 18598 10412 18604 10424
rect 18656 10412 18662 10464
rect 18782 10412 18788 10464
rect 18840 10412 18846 10464
rect 1104 10362 19136 10384
rect 1104 10310 2350 10362
rect 2402 10310 2414 10362
rect 2466 10310 2478 10362
rect 2530 10310 2542 10362
rect 2594 10310 2606 10362
rect 2658 10310 19136 10362
rect 1104 10288 19136 10310
rect 2222 10208 2228 10260
rect 2280 10248 2286 10260
rect 2409 10251 2467 10257
rect 2409 10248 2421 10251
rect 2280 10220 2421 10248
rect 2280 10208 2286 10220
rect 2409 10217 2421 10220
rect 2455 10217 2467 10251
rect 2409 10211 2467 10217
rect 15194 10208 15200 10260
rect 15252 10208 15258 10260
rect 18322 10208 18328 10260
rect 18380 10208 18386 10260
rect 842 10072 848 10124
rect 900 10112 906 10124
rect 1397 10115 1455 10121
rect 1397 10112 1409 10115
rect 900 10084 1409 10112
rect 900 10072 906 10084
rect 1397 10081 1409 10084
rect 1443 10081 1455 10115
rect 1397 10075 1455 10081
rect 1673 10115 1731 10121
rect 1673 10081 1685 10115
rect 1719 10112 1731 10115
rect 8202 10112 8208 10124
rect 1719 10084 8208 10112
rect 1719 10081 1731 10084
rect 1673 10075 1731 10081
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 16850 10072 16856 10124
rect 16908 10072 16914 10124
rect 2130 10004 2136 10056
rect 2188 10044 2194 10056
rect 2317 10047 2375 10053
rect 2317 10044 2329 10047
rect 2188 10016 2329 10044
rect 2188 10004 2194 10016
rect 2317 10013 2329 10016
rect 2363 10013 2375 10047
rect 2317 10007 2375 10013
rect 15381 10047 15439 10053
rect 15381 10013 15393 10047
rect 15427 10013 15439 10047
rect 15381 10007 15439 10013
rect 15396 9976 15424 10007
rect 15470 10004 15476 10056
rect 15528 10044 15534 10056
rect 15565 10047 15623 10053
rect 15565 10044 15577 10047
rect 15528 10016 15577 10044
rect 15528 10004 15534 10016
rect 15565 10013 15577 10016
rect 15611 10013 15623 10047
rect 15565 10007 15623 10013
rect 15657 10047 15715 10053
rect 15657 10013 15669 10047
rect 15703 10044 15715 10047
rect 15838 10044 15844 10056
rect 15703 10016 15844 10044
rect 15703 10013 15715 10016
rect 15657 10007 15715 10013
rect 15838 10004 15844 10016
rect 15896 10004 15902 10056
rect 16574 10004 16580 10056
rect 16632 10004 16638 10056
rect 18414 10004 18420 10056
rect 18472 10004 18478 10056
rect 16850 9976 16856 9988
rect 15396 9948 16856 9976
rect 16850 9936 16856 9948
rect 16908 9936 16914 9988
rect 18509 9979 18567 9985
rect 18509 9976 18521 9979
rect 18078 9948 18521 9976
rect 18509 9945 18521 9948
rect 18555 9945 18567 9979
rect 18509 9939 18567 9945
rect 1104 9818 19136 9840
rect 1104 9766 3010 9818
rect 3062 9766 3074 9818
rect 3126 9766 3138 9818
rect 3190 9766 3202 9818
rect 3254 9766 3266 9818
rect 3318 9766 19136 9818
rect 1104 9744 19136 9766
rect 1581 9707 1639 9713
rect 1581 9673 1593 9707
rect 1627 9673 1639 9707
rect 1581 9667 1639 9673
rect 1596 9636 1624 9667
rect 2133 9639 2191 9645
rect 2133 9636 2145 9639
rect 1596 9608 2145 9636
rect 2133 9605 2145 9608
rect 2179 9605 2191 9639
rect 2133 9599 2191 9605
rect 2866 9596 2872 9648
rect 2924 9596 2930 9648
rect 4154 9596 4160 9648
rect 4212 9596 4218 9648
rect 5813 9639 5871 9645
rect 5813 9636 5825 9639
rect 5382 9608 5825 9636
rect 5813 9605 5825 9608
rect 5859 9605 5871 9639
rect 5813 9599 5871 9605
rect 8110 9596 8116 9648
rect 8168 9636 8174 9648
rect 10594 9636 10600 9648
rect 8168 9608 10600 9636
rect 8168 9596 8174 9608
rect 10594 9596 10600 9608
rect 10652 9636 10658 9648
rect 12526 9636 12532 9648
rect 10652 9608 12532 9636
rect 10652 9596 10658 9608
rect 12526 9596 12532 9608
rect 12584 9636 12590 9648
rect 13173 9639 13231 9645
rect 13173 9636 13185 9639
rect 12584 9608 13185 9636
rect 12584 9596 12590 9608
rect 13173 9605 13185 9608
rect 13219 9605 13231 9639
rect 13173 9599 13231 9605
rect 17402 9596 17408 9648
rect 17460 9596 17466 9648
rect 842 9528 848 9580
rect 900 9568 906 9580
rect 1397 9571 1455 9577
rect 1397 9568 1409 9571
rect 900 9540 1409 9568
rect 900 9528 906 9540
rect 1397 9537 1409 9540
rect 1443 9537 1455 9571
rect 1397 9531 1455 9537
rect 1486 9528 1492 9580
rect 1544 9568 1550 9580
rect 1857 9571 1915 9577
rect 1857 9568 1869 9571
rect 1544 9540 1869 9568
rect 1544 9528 1550 9540
rect 1857 9537 1869 9540
rect 1903 9537 1915 9571
rect 1857 9531 1915 9537
rect 1872 9364 1900 9531
rect 5902 9528 5908 9580
rect 5960 9568 5966 9580
rect 6362 9568 6368 9580
rect 5960 9540 6368 9568
rect 5960 9528 5966 9540
rect 6362 9528 6368 9540
rect 6420 9528 6426 9580
rect 11974 9528 11980 9580
rect 12032 9528 12038 9580
rect 18693 9571 18751 9577
rect 18693 9568 18705 9571
rect 18432 9540 18705 9568
rect 3881 9503 3939 9509
rect 3881 9469 3893 9503
rect 3927 9469 3939 9503
rect 3881 9463 3939 9469
rect 3896 9432 3924 9463
rect 14182 9460 14188 9512
rect 14240 9500 14246 9512
rect 16666 9500 16672 9512
rect 14240 9472 16672 9500
rect 14240 9460 14246 9472
rect 16666 9460 16672 9472
rect 16724 9460 16730 9512
rect 16942 9460 16948 9512
rect 17000 9460 17006 9512
rect 18432 9509 18460 9540
rect 18693 9537 18705 9540
rect 18739 9537 18751 9571
rect 18693 9531 18751 9537
rect 18417 9503 18475 9509
rect 18417 9469 18429 9503
rect 18463 9469 18475 9503
rect 18417 9463 18475 9469
rect 3344 9404 3924 9432
rect 12161 9435 12219 9441
rect 2682 9364 2688 9376
rect 1872 9336 2688 9364
rect 2682 9324 2688 9336
rect 2740 9364 2746 9376
rect 3344 9364 3372 9404
rect 12161 9401 12173 9435
rect 12207 9432 12219 9435
rect 12207 9404 16574 9432
rect 12207 9401 12219 9404
rect 12161 9395 12219 9401
rect 2740 9336 3372 9364
rect 3605 9367 3663 9373
rect 2740 9324 2746 9336
rect 3605 9333 3617 9367
rect 3651 9364 3663 9367
rect 4246 9364 4252 9376
rect 3651 9336 4252 9364
rect 3651 9333 3663 9336
rect 3605 9327 3663 9333
rect 4246 9324 4252 9336
rect 4304 9324 4310 9376
rect 5626 9324 5632 9376
rect 5684 9324 5690 9376
rect 14182 9324 14188 9376
rect 14240 9364 14246 9376
rect 14461 9367 14519 9373
rect 14461 9364 14473 9367
rect 14240 9336 14473 9364
rect 14240 9324 14246 9336
rect 14461 9333 14473 9336
rect 14507 9333 14519 9367
rect 16546 9364 16574 9404
rect 17954 9364 17960 9376
rect 16546 9336 17960 9364
rect 14461 9327 14519 9333
rect 17954 9324 17960 9336
rect 18012 9324 18018 9376
rect 18322 9324 18328 9376
rect 18380 9364 18386 9376
rect 18509 9367 18567 9373
rect 18509 9364 18521 9367
rect 18380 9336 18521 9364
rect 18380 9324 18386 9336
rect 18509 9333 18521 9336
rect 18555 9333 18567 9367
rect 18509 9327 18567 9333
rect 1104 9274 19136 9296
rect 1104 9222 2350 9274
rect 2402 9222 2414 9274
rect 2466 9222 2478 9274
rect 2530 9222 2542 9274
rect 2594 9222 2606 9274
rect 2658 9222 19136 9274
rect 1104 9200 19136 9222
rect 2866 9120 2872 9172
rect 2924 9160 2930 9172
rect 2961 9163 3019 9169
rect 2961 9160 2973 9163
rect 2924 9132 2973 9160
rect 2924 9120 2930 9132
rect 2961 9129 2973 9132
rect 3007 9129 3019 9163
rect 2961 9123 3019 9129
rect 17313 9163 17371 9169
rect 17313 9129 17325 9163
rect 17359 9160 17371 9163
rect 17402 9160 17408 9172
rect 17359 9132 17408 9160
rect 17359 9129 17371 9132
rect 17313 9123 17371 9129
rect 17402 9120 17408 9132
rect 17460 9120 17466 9172
rect 18782 9120 18788 9172
rect 18840 9120 18846 9172
rect 842 9052 848 9104
rect 900 9092 906 9104
rect 1397 9095 1455 9101
rect 1397 9092 1409 9095
rect 900 9064 1409 9092
rect 900 9052 906 9064
rect 1397 9061 1409 9064
rect 1443 9061 1455 9095
rect 1397 9055 1455 9061
rect 5626 9024 5632 9036
rect 1964 8996 5632 9024
rect 1581 8959 1639 8965
rect 1581 8925 1593 8959
rect 1627 8956 1639 8959
rect 1627 8928 1808 8956
rect 1627 8925 1639 8928
rect 1581 8919 1639 8925
rect 1780 8829 1808 8928
rect 1854 8916 1860 8968
rect 1912 8956 1918 8968
rect 1964 8965 1992 8996
rect 5626 8984 5632 8996
rect 5684 8984 5690 9036
rect 8294 8984 8300 9036
rect 8352 9024 8358 9036
rect 9585 9027 9643 9033
rect 8352 8996 9352 9024
rect 8352 8984 8358 8996
rect 9324 8968 9352 8996
rect 9585 8993 9597 9027
rect 9631 9024 9643 9027
rect 9953 9027 10011 9033
rect 9953 9024 9965 9027
rect 9631 8996 9965 9024
rect 9631 8993 9643 8996
rect 9585 8987 9643 8993
rect 9953 8993 9965 8996
rect 9999 8993 10011 9027
rect 9953 8987 10011 8993
rect 1949 8959 2007 8965
rect 1949 8956 1961 8959
rect 1912 8928 1961 8956
rect 1912 8916 1918 8928
rect 1949 8925 1961 8928
rect 1995 8925 2007 8959
rect 1949 8919 2007 8925
rect 2130 8916 2136 8968
rect 2188 8956 2194 8968
rect 2869 8959 2927 8965
rect 2869 8956 2881 8959
rect 2188 8928 2881 8956
rect 2188 8916 2194 8928
rect 2869 8925 2881 8928
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 5721 8959 5779 8965
rect 5721 8925 5733 8959
rect 5767 8956 5779 8959
rect 5810 8956 5816 8968
rect 5767 8928 5816 8956
rect 5767 8925 5779 8928
rect 5721 8919 5779 8925
rect 5810 8916 5816 8928
rect 5868 8916 5874 8968
rect 8570 8916 8576 8968
rect 8628 8956 8634 8968
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8628 8928 8953 8956
rect 8628 8916 8634 8928
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 9122 8916 9128 8968
rect 9180 8916 9186 8968
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8925 9275 8959
rect 9217 8919 9275 8925
rect 9232 8888 9260 8919
rect 9306 8916 9312 8968
rect 9364 8916 9370 8968
rect 9677 8959 9735 8965
rect 9677 8925 9689 8959
rect 9723 8925 9735 8959
rect 9677 8919 9735 8925
rect 11701 8959 11759 8965
rect 11701 8925 11713 8959
rect 11747 8956 11759 8959
rect 13722 8956 13728 8968
rect 11747 8928 13728 8956
rect 11747 8925 11759 8928
rect 11701 8919 11759 8925
rect 9692 8888 9720 8919
rect 13722 8916 13728 8928
rect 13780 8916 13786 8968
rect 14182 8916 14188 8968
rect 14240 8916 14246 8968
rect 16209 8959 16267 8965
rect 16209 8925 16221 8959
rect 16255 8956 16267 8959
rect 16574 8956 16580 8968
rect 16255 8928 16580 8956
rect 16255 8925 16267 8928
rect 16209 8919 16267 8925
rect 16574 8916 16580 8928
rect 16632 8956 16638 8968
rect 17221 8959 17279 8965
rect 17221 8956 17233 8959
rect 16632 8928 17233 8956
rect 16632 8916 16638 8928
rect 17221 8925 17233 8928
rect 17267 8925 17279 8959
rect 17221 8919 17279 8925
rect 18322 8916 18328 8968
rect 18380 8916 18386 8968
rect 18598 8916 18604 8968
rect 18656 8916 18662 8968
rect 9858 8888 9864 8900
rect 9232 8860 9352 8888
rect 9692 8860 9864 8888
rect 1765 8823 1823 8829
rect 1765 8789 1777 8823
rect 1811 8789 1823 8823
rect 9324 8820 9352 8860
rect 9858 8848 9864 8860
rect 9916 8848 9922 8900
rect 11609 8891 11667 8897
rect 11609 8888 11621 8891
rect 11178 8860 11621 8888
rect 11609 8857 11621 8860
rect 11655 8857 11667 8891
rect 11609 8851 11667 8857
rect 14461 8891 14519 8897
rect 14461 8857 14473 8891
rect 14507 8857 14519 8891
rect 16117 8891 16175 8897
rect 16117 8888 16129 8891
rect 15686 8860 16129 8888
rect 14461 8851 14519 8857
rect 16117 8857 16129 8860
rect 16163 8857 16175 8891
rect 16117 8851 16175 8857
rect 9674 8820 9680 8832
rect 9324 8792 9680 8820
rect 1765 8783 1823 8789
rect 9674 8780 9680 8792
rect 9732 8780 9738 8832
rect 9766 8780 9772 8832
rect 9824 8820 9830 8832
rect 11425 8823 11483 8829
rect 11425 8820 11437 8823
rect 9824 8792 11437 8820
rect 9824 8780 9830 8792
rect 11425 8789 11437 8792
rect 11471 8820 11483 8823
rect 11974 8820 11980 8832
rect 11471 8792 11980 8820
rect 11471 8789 11483 8792
rect 11425 8783 11483 8789
rect 11974 8780 11980 8792
rect 12032 8780 12038 8832
rect 14476 8820 14504 8851
rect 15378 8820 15384 8832
rect 14476 8792 15384 8820
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 15933 8823 15991 8829
rect 15933 8789 15945 8823
rect 15979 8820 15991 8823
rect 16022 8820 16028 8832
rect 15979 8792 16028 8820
rect 15979 8789 15991 8792
rect 15933 8783 15991 8789
rect 16022 8780 16028 8792
rect 16080 8780 16086 8832
rect 18506 8780 18512 8832
rect 18564 8780 18570 8832
rect 1104 8730 19136 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 19136 8730
rect 1104 8656 19136 8678
rect 2682 8576 2688 8628
rect 2740 8576 2746 8628
rect 4157 8619 4215 8625
rect 4157 8585 4169 8619
rect 4203 8616 4215 8619
rect 4525 8619 4583 8625
rect 4525 8616 4537 8619
rect 4203 8588 4537 8616
rect 4203 8585 4215 8588
rect 4157 8579 4215 8585
rect 4525 8585 4537 8588
rect 4571 8585 4583 8619
rect 4525 8579 4583 8585
rect 9122 8576 9128 8628
rect 9180 8616 9186 8628
rect 9401 8619 9459 8625
rect 9401 8616 9413 8619
rect 9180 8588 9413 8616
rect 9180 8576 9186 8588
rect 9401 8585 9413 8588
rect 9447 8585 9459 8619
rect 9401 8579 9459 8585
rect 2222 8508 2228 8560
rect 2280 8508 2286 8560
rect 2700 8548 2728 8576
rect 5810 8548 5816 8560
rect 2700 8520 5816 8548
rect 3160 8489 3188 8520
rect 5810 8508 5816 8520
rect 5868 8548 5874 8560
rect 6365 8551 6423 8557
rect 6365 8548 6377 8551
rect 5868 8520 6377 8548
rect 5868 8508 5874 8520
rect 6365 8517 6377 8520
rect 6411 8517 6423 8551
rect 6365 8511 6423 8517
rect 16209 8551 16267 8557
rect 16209 8517 16221 8551
rect 16255 8548 16267 8551
rect 17402 8548 17408 8560
rect 16255 8520 17408 8548
rect 16255 8517 16267 8520
rect 16209 8511 16267 8517
rect 17402 8508 17408 8520
rect 17460 8508 17466 8560
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8449 3203 8483
rect 3145 8443 3203 8449
rect 4246 8440 4252 8492
rect 4304 8440 4310 8492
rect 4614 8440 4620 8492
rect 4672 8440 4678 8492
rect 8110 8440 8116 8492
rect 8168 8440 8174 8492
rect 9306 8440 9312 8492
rect 9364 8480 9370 8492
rect 9615 8483 9673 8489
rect 9615 8480 9627 8483
rect 9364 8452 9627 8480
rect 9364 8440 9370 8452
rect 9615 8449 9627 8452
rect 9661 8449 9673 8483
rect 9615 8443 9673 8449
rect 9766 8440 9772 8492
rect 9824 8440 9830 8492
rect 9858 8440 9864 8492
rect 9916 8480 9922 8492
rect 13173 8483 13231 8489
rect 13173 8480 13185 8483
rect 9916 8452 13185 8480
rect 9916 8440 9922 8452
rect 13173 8449 13185 8452
rect 13219 8480 13231 8483
rect 14182 8480 14188 8492
rect 13219 8452 14188 8480
rect 13219 8449 13231 8452
rect 13173 8443 13231 8449
rect 14182 8440 14188 8452
rect 14240 8440 14246 8492
rect 16666 8440 16672 8492
rect 16724 8480 16730 8492
rect 16853 8483 16911 8489
rect 16853 8480 16865 8483
rect 16724 8452 16865 8480
rect 16724 8440 16730 8452
rect 16853 8449 16865 8452
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 18230 8440 18236 8492
rect 18288 8440 18294 8492
rect 2866 8372 2872 8424
rect 2924 8372 2930 8424
rect 3789 8415 3847 8421
rect 3789 8381 3801 8415
rect 3835 8412 3847 8415
rect 15565 8415 15623 8421
rect 3835 8384 4292 8412
rect 3835 8381 3847 8384
rect 3789 8375 3847 8381
rect 4264 8356 4292 8384
rect 15565 8381 15577 8415
rect 15611 8412 15623 8415
rect 15654 8412 15660 8424
rect 15611 8384 15660 8412
rect 15611 8381 15623 8384
rect 15565 8375 15623 8381
rect 15654 8372 15660 8384
rect 15712 8372 15718 8424
rect 15746 8372 15752 8424
rect 15804 8372 15810 8424
rect 17126 8372 17132 8424
rect 17184 8372 17190 8424
rect 3973 8347 4031 8353
rect 3973 8313 3985 8347
rect 4019 8344 4031 8347
rect 4154 8344 4160 8356
rect 4019 8316 4160 8344
rect 4019 8313 4031 8316
rect 3973 8307 4031 8313
rect 4154 8304 4160 8316
rect 4212 8304 4218 8356
rect 4246 8304 4252 8356
rect 4304 8304 4310 8356
rect 1397 8279 1455 8285
rect 1397 8245 1409 8279
rect 1443 8276 1455 8279
rect 1762 8276 1768 8288
rect 1443 8248 1768 8276
rect 1443 8245 1455 8248
rect 1397 8239 1455 8245
rect 1762 8236 1768 8248
rect 1820 8236 1826 8288
rect 18138 8236 18144 8288
rect 18196 8276 18202 8288
rect 18601 8279 18659 8285
rect 18601 8276 18613 8279
rect 18196 8248 18613 8276
rect 18196 8236 18202 8248
rect 18601 8245 18613 8248
rect 18647 8245 18659 8279
rect 18601 8239 18659 8245
rect 1104 8186 19136 8208
rect 1104 8134 2350 8186
rect 2402 8134 2414 8186
rect 2466 8134 2478 8186
rect 2530 8134 2542 8186
rect 2594 8134 2606 8186
rect 2658 8134 19136 8186
rect 1104 8112 19136 8134
rect 1302 8032 1308 8084
rect 1360 8072 1366 8084
rect 1397 8075 1455 8081
rect 1397 8072 1409 8075
rect 1360 8044 1409 8072
rect 1360 8032 1366 8044
rect 1397 8041 1409 8044
rect 1443 8041 1455 8075
rect 1397 8035 1455 8041
rect 2222 8032 2228 8084
rect 2280 8072 2286 8084
rect 2317 8075 2375 8081
rect 2317 8072 2329 8075
rect 2280 8044 2329 8072
rect 2280 8032 2286 8044
rect 2317 8041 2329 8044
rect 2363 8041 2375 8075
rect 8570 8072 8576 8084
rect 2317 8035 2375 8041
rect 3804 8044 8576 8072
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7868 1639 7871
rect 1673 7871 1731 7877
rect 1673 7868 1685 7871
rect 1627 7840 1685 7868
rect 1627 7837 1639 7840
rect 1581 7831 1639 7837
rect 1673 7837 1685 7840
rect 1719 7837 1731 7871
rect 1673 7831 1731 7837
rect 1762 7828 1768 7880
rect 1820 7868 1826 7880
rect 2041 7871 2099 7877
rect 2041 7868 2053 7871
rect 1820 7840 2053 7868
rect 1820 7828 1826 7840
rect 2041 7837 2053 7840
rect 2087 7837 2099 7871
rect 2041 7831 2099 7837
rect 1854 7760 1860 7812
rect 1912 7760 1918 7812
rect 2056 7800 2084 7831
rect 2130 7828 2136 7880
rect 2188 7868 2194 7880
rect 2409 7871 2467 7877
rect 2409 7868 2421 7871
rect 2188 7840 2421 7868
rect 2188 7828 2194 7840
rect 2409 7837 2421 7840
rect 2455 7868 2467 7871
rect 2590 7868 2596 7880
rect 2455 7840 2596 7868
rect 2455 7837 2467 7840
rect 2409 7831 2467 7837
rect 2590 7828 2596 7840
rect 2648 7828 2654 7880
rect 2685 7871 2743 7877
rect 2685 7837 2697 7871
rect 2731 7837 2743 7871
rect 2685 7831 2743 7837
rect 2700 7800 2728 7831
rect 3602 7828 3608 7880
rect 3660 7868 3666 7880
rect 3804 7877 3832 8044
rect 8570 8032 8576 8044
rect 8628 8032 8634 8084
rect 15746 8032 15752 8084
rect 15804 8072 15810 8084
rect 16117 8075 16175 8081
rect 16117 8072 16129 8075
rect 15804 8044 16129 8072
rect 15804 8032 15810 8044
rect 16117 8041 16129 8044
rect 16163 8041 16175 8075
rect 16117 8035 16175 8041
rect 17037 8075 17095 8081
rect 17037 8041 17049 8075
rect 17083 8072 17095 8075
rect 17126 8072 17132 8084
rect 17083 8044 17132 8072
rect 17083 8041 17095 8044
rect 17037 8035 17095 8041
rect 17126 8032 17132 8044
rect 17184 8032 17190 8084
rect 18230 8032 18236 8084
rect 18288 8072 18294 8084
rect 18325 8075 18383 8081
rect 18325 8072 18337 8075
rect 18288 8044 18337 8072
rect 18288 8032 18294 8044
rect 18325 8041 18337 8044
rect 18371 8041 18383 8075
rect 18325 8035 18383 8041
rect 4154 7964 4160 8016
rect 4212 7964 4218 8016
rect 3878 7896 3884 7948
rect 3936 7896 3942 7948
rect 3970 7896 3976 7948
rect 4028 7896 4034 7948
rect 4249 7939 4307 7945
rect 4249 7905 4261 7939
rect 4295 7936 4307 7939
rect 5810 7936 5816 7948
rect 4295 7908 5816 7936
rect 4295 7905 4307 7908
rect 4249 7899 4307 7905
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 14090 7896 14096 7948
rect 14148 7896 14154 7948
rect 15378 7896 15384 7948
rect 15436 7936 15442 7948
rect 15436 7908 17816 7936
rect 15436 7896 15442 7908
rect 3789 7871 3847 7877
rect 3789 7868 3801 7871
rect 3660 7840 3801 7868
rect 3660 7828 3666 7840
rect 3789 7837 3801 7840
rect 3835 7837 3847 7871
rect 3789 7831 3847 7837
rect 6822 7828 6828 7880
rect 6880 7868 6886 7880
rect 9122 7868 9128 7880
rect 6880 7840 9128 7868
rect 6880 7828 6886 7840
rect 9122 7828 9128 7840
rect 9180 7828 9186 7880
rect 13446 7828 13452 7880
rect 13504 7868 13510 7880
rect 13722 7868 13728 7880
rect 13504 7840 13728 7868
rect 13504 7828 13510 7840
rect 13722 7828 13728 7840
rect 13780 7828 13786 7880
rect 15930 7828 15936 7880
rect 15988 7828 15994 7880
rect 16022 7828 16028 7880
rect 16080 7868 16086 7880
rect 17328 7877 17356 7908
rect 17313 7871 17371 7877
rect 16080 7840 16125 7868
rect 16080 7828 16086 7840
rect 17313 7837 17325 7871
rect 17359 7837 17371 7871
rect 17313 7831 17371 7837
rect 17402 7828 17408 7880
rect 17460 7828 17466 7880
rect 17497 7871 17555 7877
rect 17497 7837 17509 7871
rect 17543 7837 17555 7871
rect 17497 7831 17555 7837
rect 2056 7772 2728 7800
rect 4087 7803 4145 7809
rect 4087 7769 4099 7803
rect 4133 7800 4145 7803
rect 4525 7803 4583 7809
rect 4525 7800 4537 7803
rect 4133 7772 4537 7800
rect 4133 7769 4145 7772
rect 4087 7763 4145 7769
rect 4525 7769 4537 7772
rect 4571 7769 4583 7803
rect 4525 7763 4583 7769
rect 5534 7760 5540 7812
rect 5592 7760 5598 7812
rect 14369 7803 14427 7809
rect 14369 7769 14381 7803
rect 14415 7800 14427 7803
rect 14642 7800 14648 7812
rect 14415 7772 14648 7800
rect 14415 7769 14427 7772
rect 14369 7763 14427 7769
rect 14642 7760 14648 7772
rect 14700 7760 14706 7812
rect 17512 7800 17540 7831
rect 17678 7828 17684 7880
rect 17736 7828 17742 7880
rect 17788 7868 17816 7908
rect 18046 7868 18052 7880
rect 17788 7840 18052 7868
rect 18046 7828 18052 7840
rect 18104 7828 18110 7880
rect 18138 7828 18144 7880
rect 18196 7828 18202 7880
rect 18417 7871 18475 7877
rect 18417 7837 18429 7871
rect 18463 7837 18475 7871
rect 18417 7831 18475 7837
rect 17773 7803 17831 7809
rect 17773 7800 17785 7803
rect 14752 7772 14858 7800
rect 17512 7772 17785 7800
rect 2498 7692 2504 7744
rect 2556 7692 2562 7744
rect 4798 7692 4804 7744
rect 4856 7732 4862 7744
rect 5997 7735 6055 7741
rect 5997 7732 6009 7735
rect 4856 7704 6009 7732
rect 4856 7692 4862 7704
rect 5997 7701 6009 7704
rect 6043 7701 6055 7735
rect 5997 7695 6055 7701
rect 9030 7692 9036 7744
rect 9088 7692 9094 7744
rect 13817 7735 13875 7741
rect 13817 7701 13829 7735
rect 13863 7732 13875 7735
rect 14752 7732 14780 7772
rect 17773 7769 17785 7772
rect 17819 7769 17831 7803
rect 17773 7763 17831 7769
rect 13863 7704 14780 7732
rect 13863 7701 13875 7704
rect 13817 7695 13875 7701
rect 15746 7692 15752 7744
rect 15804 7732 15810 7744
rect 15841 7735 15899 7741
rect 15841 7732 15853 7735
rect 15804 7704 15853 7732
rect 15804 7692 15810 7704
rect 15841 7701 15853 7704
rect 15887 7701 15899 7735
rect 15841 7695 15899 7701
rect 16574 7692 16580 7744
rect 16632 7732 16638 7744
rect 18432 7732 18460 7831
rect 18598 7828 18604 7880
rect 18656 7828 18662 7880
rect 16632 7704 18460 7732
rect 16632 7692 16638 7704
rect 18782 7692 18788 7744
rect 18840 7692 18846 7744
rect 1104 7642 19136 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 19136 7642
rect 1104 7568 19136 7590
rect 1302 7488 1308 7540
rect 1360 7528 1366 7540
rect 1397 7531 1455 7537
rect 1397 7528 1409 7531
rect 1360 7500 1409 7528
rect 1360 7488 1366 7500
rect 1397 7497 1409 7500
rect 1443 7497 1455 7531
rect 1397 7491 1455 7497
rect 2866 7488 2872 7540
rect 2924 7528 2930 7540
rect 3329 7531 3387 7537
rect 3329 7528 3341 7531
rect 2924 7500 3341 7528
rect 2924 7488 2930 7500
rect 3329 7497 3341 7500
rect 3375 7497 3387 7531
rect 3329 7491 3387 7497
rect 3878 7488 3884 7540
rect 3936 7528 3942 7540
rect 4709 7531 4767 7537
rect 4709 7528 4721 7531
rect 3936 7500 4721 7528
rect 3936 7488 3942 7500
rect 4709 7497 4721 7500
rect 4755 7497 4767 7531
rect 4709 7491 4767 7497
rect 5445 7531 5503 7537
rect 5445 7497 5457 7531
rect 5491 7528 5503 7531
rect 5534 7528 5540 7540
rect 5491 7500 5540 7528
rect 5491 7497 5503 7500
rect 5445 7491 5503 7497
rect 5534 7488 5540 7500
rect 5592 7488 5598 7540
rect 5902 7488 5908 7540
rect 5960 7528 5966 7540
rect 6822 7528 6828 7540
rect 5960 7500 6828 7528
rect 5960 7488 5966 7500
rect 6822 7488 6828 7500
rect 6880 7528 6886 7540
rect 6880 7500 7420 7528
rect 6880 7488 6886 7500
rect 4433 7463 4491 7469
rect 4433 7429 4445 7463
rect 4479 7460 4491 7463
rect 4614 7460 4620 7472
rect 4479 7432 4620 7460
rect 4479 7429 4491 7432
rect 4433 7423 4491 7429
rect 4614 7420 4620 7432
rect 4672 7460 4678 7472
rect 4672 7432 6868 7460
rect 4672 7420 4678 7432
rect 1581 7395 1639 7401
rect 1581 7361 1593 7395
rect 1627 7392 1639 7395
rect 2498 7392 2504 7404
rect 1627 7364 2504 7392
rect 1627 7361 1639 7364
rect 1581 7355 1639 7361
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7361 3663 7395
rect 3605 7355 3663 7361
rect 3620 7324 3648 7355
rect 3694 7352 3700 7404
rect 3752 7352 3758 7404
rect 3789 7395 3847 7401
rect 3789 7361 3801 7395
rect 3835 7392 3847 7395
rect 3878 7392 3884 7404
rect 3835 7364 3884 7392
rect 3835 7361 3847 7364
rect 3789 7355 3847 7361
rect 3878 7352 3884 7364
rect 3936 7352 3942 7404
rect 3973 7395 4031 7401
rect 3973 7361 3985 7395
rect 4019 7361 4031 7395
rect 3973 7355 4031 7361
rect 3988 7324 4016 7355
rect 4246 7352 4252 7404
rect 4304 7352 4310 7404
rect 4522 7352 4528 7404
rect 4580 7352 4586 7404
rect 4798 7352 4804 7404
rect 4856 7352 4862 7404
rect 5537 7395 5595 7401
rect 5537 7361 5549 7395
rect 5583 7392 5595 7395
rect 5902 7392 5908 7404
rect 5583 7364 5908 7392
rect 5583 7361 5595 7364
rect 5537 7355 5595 7361
rect 5902 7352 5908 7364
rect 5960 7352 5966 7404
rect 6840 7401 6868 7432
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7361 6791 7395
rect 6733 7355 6791 7361
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7392 6883 7395
rect 7282 7392 7288 7404
rect 6871 7364 7288 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 4816 7324 4844 7352
rect 3620 7296 3832 7324
rect 3988 7296 4844 7324
rect 3804 7268 3832 7296
rect 3786 7216 3792 7268
rect 3844 7216 3850 7268
rect 4246 7216 4252 7268
rect 4304 7256 4310 7268
rect 5994 7256 6000 7268
rect 4304 7228 6000 7256
rect 4304 7216 4310 7228
rect 5994 7216 6000 7228
rect 6052 7256 6058 7268
rect 6748 7256 6776 7355
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 7392 7401 7420 7500
rect 14642 7488 14648 7540
rect 14700 7488 14706 7540
rect 15013 7531 15071 7537
rect 15013 7497 15025 7531
rect 15059 7528 15071 7531
rect 15197 7531 15255 7537
rect 15197 7528 15209 7531
rect 15059 7500 15209 7528
rect 15059 7497 15071 7500
rect 15013 7491 15071 7497
rect 15197 7497 15209 7500
rect 15243 7497 15255 7531
rect 15197 7491 15255 7497
rect 15286 7488 15292 7540
rect 15344 7528 15350 7540
rect 17678 7528 17684 7540
rect 15344 7500 17684 7528
rect 15344 7488 15350 7500
rect 17678 7488 17684 7500
rect 17736 7488 17742 7540
rect 8021 7463 8079 7469
rect 8021 7429 8033 7463
rect 8067 7460 8079 7463
rect 8294 7460 8300 7472
rect 8067 7432 8300 7460
rect 8067 7429 8079 7432
rect 8021 7423 8079 7429
rect 8294 7420 8300 7432
rect 8352 7420 8358 7472
rect 9030 7420 9036 7472
rect 9088 7420 9094 7472
rect 15746 7460 15752 7472
rect 15120 7432 15752 7460
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 12897 7395 12955 7401
rect 12897 7361 12909 7395
rect 12943 7392 12955 7395
rect 13722 7392 13728 7404
rect 12943 7364 13728 7392
rect 12943 7361 12955 7364
rect 12897 7355 12955 7361
rect 13722 7352 13728 7364
rect 13780 7352 13786 7404
rect 15120 7401 15148 7432
rect 15746 7420 15752 7432
rect 15804 7420 15810 7472
rect 15841 7463 15899 7469
rect 15841 7429 15853 7463
rect 15887 7460 15899 7463
rect 17402 7460 17408 7472
rect 15887 7432 17408 7460
rect 15887 7429 15899 7432
rect 15841 7423 15899 7429
rect 17402 7420 17408 7432
rect 17460 7420 17466 7472
rect 14829 7395 14887 7401
rect 14829 7361 14841 7395
rect 14875 7361 14887 7395
rect 14829 7355 14887 7361
rect 15105 7395 15163 7401
rect 15105 7361 15117 7395
rect 15151 7361 15163 7395
rect 15105 7355 15163 7361
rect 15197 7395 15255 7401
rect 15197 7361 15209 7395
rect 15243 7392 15255 7395
rect 15286 7392 15292 7404
rect 15243 7364 15292 7392
rect 15243 7361 15255 7364
rect 15197 7355 15255 7361
rect 6917 7327 6975 7333
rect 6917 7324 6929 7327
rect 6840 7296 6929 7324
rect 6840 7268 6868 7296
rect 6917 7293 6929 7296
rect 6963 7293 6975 7327
rect 6917 7287 6975 7293
rect 7558 7284 7564 7336
rect 7616 7324 7622 7336
rect 7745 7327 7803 7333
rect 7745 7324 7757 7327
rect 7616 7296 7757 7324
rect 7616 7284 7622 7296
rect 7745 7293 7757 7296
rect 7791 7293 7803 7327
rect 7745 7287 7803 7293
rect 9582 7284 9588 7336
rect 9640 7284 9646 7336
rect 9766 7284 9772 7336
rect 9824 7284 9830 7336
rect 14844 7324 14872 7355
rect 15286 7352 15292 7364
rect 15344 7352 15350 7404
rect 15378 7352 15384 7404
rect 15436 7352 15442 7404
rect 15470 7352 15476 7404
rect 15528 7392 15534 7404
rect 16022 7392 16028 7404
rect 15528 7364 16028 7392
rect 15528 7352 15534 7364
rect 16022 7352 16028 7364
rect 16080 7352 16086 7404
rect 18138 7352 18144 7404
rect 18196 7352 18202 7404
rect 18322 7352 18328 7404
rect 18380 7392 18386 7404
rect 18601 7395 18659 7401
rect 18601 7392 18613 7395
rect 18380 7364 18613 7392
rect 18380 7352 18386 7364
rect 18601 7361 18613 7364
rect 18647 7361 18659 7395
rect 18601 7355 18659 7361
rect 15838 7324 15844 7336
rect 14844 7296 15844 7324
rect 15838 7284 15844 7296
rect 15896 7324 15902 7336
rect 15896 7296 16068 7324
rect 15896 7284 15902 7296
rect 6052 7228 6776 7256
rect 6052 7216 6058 7228
rect 6822 7216 6828 7268
rect 6880 7216 6886 7268
rect 16040 7265 16068 7296
rect 16025 7259 16083 7265
rect 16025 7225 16037 7259
rect 16071 7225 16083 7259
rect 16025 7219 16083 7225
rect 4062 7148 4068 7200
rect 4120 7148 4126 7200
rect 6362 7148 6368 7200
rect 6420 7148 6426 7200
rect 7098 7148 7104 7200
rect 7156 7188 7162 7200
rect 7285 7191 7343 7197
rect 7285 7188 7297 7191
rect 7156 7160 7297 7188
rect 7156 7148 7162 7160
rect 7285 7157 7297 7160
rect 7331 7157 7343 7191
rect 7285 7151 7343 7157
rect 9490 7148 9496 7200
rect 9548 7148 9554 7200
rect 9674 7148 9680 7200
rect 9732 7188 9738 7200
rect 9953 7191 10011 7197
rect 9953 7188 9965 7191
rect 9732 7160 9965 7188
rect 9732 7148 9738 7160
rect 9953 7157 9965 7160
rect 9999 7157 10011 7191
rect 9953 7151 10011 7157
rect 15378 7148 15384 7200
rect 15436 7188 15442 7200
rect 15841 7191 15899 7197
rect 15841 7188 15853 7191
rect 15436 7160 15853 7188
rect 15436 7148 15442 7160
rect 15841 7157 15853 7160
rect 15887 7157 15899 7191
rect 15841 7151 15899 7157
rect 18325 7191 18383 7197
rect 18325 7157 18337 7191
rect 18371 7188 18383 7191
rect 18506 7188 18512 7200
rect 18371 7160 18512 7188
rect 18371 7157 18383 7160
rect 18325 7151 18383 7157
rect 18506 7148 18512 7160
rect 18564 7148 18570 7200
rect 18782 7148 18788 7200
rect 18840 7148 18846 7200
rect 1104 7098 19136 7120
rect 1104 7046 2350 7098
rect 2402 7046 2414 7098
rect 2466 7046 2478 7098
rect 2530 7046 2542 7098
rect 2594 7046 2606 7098
rect 2658 7046 19136 7098
rect 1104 7024 19136 7046
rect 3970 6944 3976 6996
rect 4028 6944 4034 6996
rect 5800 6987 5858 6993
rect 5800 6953 5812 6987
rect 5846 6984 5858 6987
rect 6362 6984 6368 6996
rect 5846 6956 6368 6984
rect 5846 6953 5858 6956
rect 5800 6947 5858 6953
rect 6362 6944 6368 6956
rect 6420 6944 6426 6996
rect 7282 6944 7288 6996
rect 7340 6944 7346 6996
rect 15838 6993 15844 6996
rect 12424 6987 12482 6993
rect 12424 6953 12436 6987
rect 12470 6984 12482 6987
rect 14093 6987 14151 6993
rect 14093 6984 14105 6987
rect 12470 6956 14105 6984
rect 12470 6953 12482 6956
rect 12424 6947 12482 6953
rect 14093 6953 14105 6956
rect 14139 6953 14151 6987
rect 14093 6947 14151 6953
rect 15828 6987 15844 6993
rect 15828 6953 15840 6987
rect 15828 6947 15844 6953
rect 15838 6944 15844 6947
rect 15896 6944 15902 6996
rect 18322 6944 18328 6996
rect 18380 6944 18386 6996
rect 18598 6944 18604 6996
rect 18656 6944 18662 6996
rect 9401 6919 9459 6925
rect 9401 6885 9413 6919
rect 9447 6916 9459 6919
rect 9766 6916 9772 6928
rect 9447 6888 9772 6916
rect 9447 6885 9459 6888
rect 9401 6879 9459 6885
rect 9766 6876 9772 6888
rect 9824 6876 9830 6928
rect 3694 6808 3700 6860
rect 3752 6848 3758 6860
rect 3752 6820 3924 6848
rect 3752 6808 3758 6820
rect 3896 6792 3924 6820
rect 4062 6808 4068 6860
rect 4120 6808 4126 6860
rect 5537 6851 5595 6857
rect 5537 6817 5549 6851
rect 5583 6848 5595 6851
rect 5810 6848 5816 6860
rect 5583 6820 5816 6848
rect 5583 6817 5595 6820
rect 5537 6811 5595 6817
rect 5810 6808 5816 6820
rect 5868 6808 5874 6860
rect 12161 6851 12219 6857
rect 12161 6817 12173 6851
rect 12207 6848 12219 6851
rect 14090 6848 14096 6860
rect 12207 6820 14096 6848
rect 12207 6817 12219 6820
rect 12161 6811 12219 6817
rect 14090 6808 14096 6820
rect 14148 6808 14154 6860
rect 14737 6851 14795 6857
rect 14737 6848 14749 6851
rect 14200 6820 14749 6848
rect 1394 6740 1400 6792
rect 1452 6740 1458 6792
rect 3786 6740 3792 6792
rect 3844 6740 3850 6792
rect 3878 6740 3884 6792
rect 3936 6740 3942 6792
rect 3970 6740 3976 6792
rect 4028 6780 4034 6792
rect 4157 6783 4215 6789
rect 4157 6780 4169 6783
rect 4028 6752 4169 6780
rect 4028 6740 4034 6752
rect 4157 6749 4169 6752
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 8294 6740 8300 6792
rect 8352 6780 8358 6792
rect 8389 6783 8447 6789
rect 8389 6780 8401 6783
rect 8352 6752 8401 6780
rect 8352 6740 8358 6752
rect 8389 6749 8401 6752
rect 8435 6749 8447 6783
rect 8389 6743 8447 6749
rect 8570 6740 8576 6792
rect 8628 6740 8634 6792
rect 9030 6740 9036 6792
rect 9088 6740 9094 6792
rect 9187 6783 9245 6789
rect 9187 6749 9199 6783
rect 9233 6780 9245 6783
rect 9490 6780 9496 6792
rect 9233 6752 9496 6780
rect 9233 6749 9245 6752
rect 9187 6743 9245 6749
rect 9490 6740 9496 6752
rect 9548 6740 9554 6792
rect 14200 6780 14228 6820
rect 14737 6817 14749 6820
rect 14783 6817 14795 6851
rect 16574 6848 16580 6860
rect 14737 6811 14795 6817
rect 14844 6820 16580 6848
rect 13570 6752 14228 6780
rect 14277 6783 14335 6789
rect 14277 6749 14289 6783
rect 14323 6780 14335 6783
rect 14366 6780 14372 6792
rect 14323 6752 14372 6780
rect 14323 6749 14335 6752
rect 14277 6743 14335 6749
rect 14366 6740 14372 6752
rect 14424 6740 14430 6792
rect 14553 6783 14611 6789
rect 14553 6758 14565 6783
rect 14476 6749 14565 6758
rect 14599 6780 14611 6783
rect 14642 6780 14648 6792
rect 14599 6752 14648 6780
rect 14599 6749 14611 6752
rect 14476 6743 14611 6749
rect 14476 6730 14596 6743
rect 14642 6740 14648 6752
rect 14700 6740 14706 6792
rect 14844 6789 14872 6820
rect 16574 6808 16580 6820
rect 16632 6848 16638 6860
rect 17218 6848 17224 6860
rect 16632 6820 17224 6848
rect 16632 6808 16638 6820
rect 17218 6808 17224 6820
rect 17276 6808 17282 6860
rect 17313 6851 17371 6857
rect 17313 6817 17325 6851
rect 17359 6848 17371 6851
rect 17359 6820 18184 6848
rect 17359 6817 17371 6820
rect 17313 6811 17371 6817
rect 14829 6783 14887 6789
rect 14829 6749 14841 6783
rect 14875 6749 14887 6783
rect 14829 6743 14887 6749
rect 15562 6740 15568 6792
rect 15620 6740 15626 6792
rect 18156 6789 18184 6820
rect 18141 6783 18199 6789
rect 18141 6749 18153 6783
rect 18187 6749 18199 6783
rect 18141 6743 18199 6749
rect 18417 6783 18475 6789
rect 18417 6749 18429 6783
rect 18463 6780 18475 6783
rect 18598 6780 18604 6792
rect 18463 6752 18604 6780
rect 18463 6749 18475 6752
rect 18417 6743 18475 6749
rect 18598 6740 18604 6752
rect 18656 6740 18662 6792
rect 1670 6672 1676 6724
rect 1728 6672 1734 6724
rect 2406 6672 2412 6724
rect 2464 6672 2470 6724
rect 7098 6712 7104 6724
rect 7038 6684 7104 6712
rect 7098 6672 7104 6684
rect 7156 6672 7162 6724
rect 14476 6712 14504 6730
rect 13924 6684 14504 6712
rect 3145 6647 3203 6653
rect 3145 6613 3157 6647
rect 3191 6644 3203 6647
rect 3418 6644 3424 6656
rect 3191 6616 3424 6644
rect 3191 6613 3203 6616
rect 3145 6607 3203 6613
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 8573 6647 8631 6653
rect 8573 6613 8585 6647
rect 8619 6644 8631 6647
rect 9306 6644 9312 6656
rect 8619 6616 9312 6644
rect 8619 6613 8631 6616
rect 8573 6607 8631 6613
rect 9306 6604 9312 6616
rect 9364 6604 9370 6656
rect 13924 6653 13952 6684
rect 16850 6672 16856 6724
rect 16908 6672 16914 6724
rect 13909 6647 13967 6653
rect 13909 6613 13921 6647
rect 13955 6613 13967 6647
rect 13909 6607 13967 6613
rect 14458 6604 14464 6656
rect 14516 6604 14522 6656
rect 1104 6554 19136 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 19136 6554
rect 1104 6480 19136 6502
rect 2406 6400 2412 6452
rect 2464 6400 2470 6452
rect 3421 6443 3479 6449
rect 3421 6409 3433 6443
rect 3467 6440 3479 6443
rect 3970 6440 3976 6452
rect 3467 6412 3976 6440
rect 3467 6409 3479 6412
rect 3421 6403 3479 6409
rect 3970 6400 3976 6412
rect 4028 6400 4034 6452
rect 9309 6443 9367 6449
rect 9309 6409 9321 6443
rect 9355 6440 9367 6443
rect 9582 6440 9588 6452
rect 9355 6412 9588 6440
rect 9355 6409 9367 6412
rect 9309 6403 9367 6409
rect 9582 6400 9588 6412
rect 9640 6400 9646 6452
rect 14458 6400 14464 6452
rect 14516 6400 14522 6452
rect 14550 6400 14556 6452
rect 14608 6440 14614 6452
rect 16761 6443 16819 6449
rect 14608 6412 16574 6440
rect 14608 6400 14614 6412
rect 16546 6384 16574 6412
rect 16761 6409 16773 6443
rect 16807 6440 16819 6443
rect 16850 6440 16856 6452
rect 16807 6412 16856 6440
rect 16807 6409 16819 6412
rect 16761 6403 16819 6409
rect 16850 6400 16856 6412
rect 16908 6400 16914 6452
rect 18046 6400 18052 6452
rect 18104 6440 18110 6452
rect 18601 6443 18659 6449
rect 18601 6440 18613 6443
rect 18104 6412 18613 6440
rect 18104 6400 18110 6412
rect 18601 6409 18613 6412
rect 18647 6409 18659 6443
rect 18601 6403 18659 6409
rect 9493 6375 9551 6381
rect 9493 6372 9505 6375
rect 9062 6344 9505 6372
rect 9493 6341 9505 6344
rect 9539 6341 9551 6375
rect 9493 6335 9551 6341
rect 12526 6332 12532 6384
rect 12584 6332 12590 6384
rect 15286 6372 15292 6384
rect 14384 6344 15292 6372
rect 842 6264 848 6316
rect 900 6304 906 6316
rect 1489 6307 1547 6313
rect 1489 6304 1501 6307
rect 900 6276 1501 6304
rect 900 6264 906 6276
rect 1489 6273 1501 6276
rect 1535 6273 1547 6307
rect 1489 6267 1547 6273
rect 1578 6264 1584 6316
rect 1636 6304 1642 6316
rect 1765 6307 1823 6313
rect 1765 6304 1777 6307
rect 1636 6276 1777 6304
rect 1636 6264 1642 6276
rect 1765 6273 1777 6276
rect 1811 6273 1823 6307
rect 1765 6267 1823 6273
rect 2130 6264 2136 6316
rect 2188 6304 2194 6316
rect 2317 6307 2375 6313
rect 2317 6304 2329 6307
rect 2188 6276 2329 6304
rect 2188 6264 2194 6276
rect 2317 6273 2329 6276
rect 2363 6304 2375 6307
rect 2682 6304 2688 6316
rect 2363 6276 2688 6304
rect 2363 6273 2375 6276
rect 2317 6267 2375 6273
rect 2682 6264 2688 6276
rect 2740 6264 2746 6316
rect 2774 6264 2780 6316
rect 2832 6304 2838 6316
rect 2961 6307 3019 6313
rect 2961 6304 2973 6307
rect 2832 6276 2973 6304
rect 2832 6264 2838 6276
rect 2961 6273 2973 6276
rect 3007 6304 3019 6307
rect 3694 6304 3700 6316
rect 3007 6276 3700 6304
rect 3007 6273 3019 6276
rect 2961 6267 3019 6273
rect 3694 6264 3700 6276
rect 3752 6264 3758 6316
rect 9122 6264 9128 6316
rect 9180 6304 9186 6316
rect 9585 6307 9643 6313
rect 9585 6304 9597 6307
rect 9180 6276 9597 6304
rect 9180 6264 9186 6276
rect 9585 6273 9597 6276
rect 9631 6304 9643 6307
rect 9766 6304 9772 6316
rect 9631 6276 9772 6304
rect 9631 6273 9643 6276
rect 9585 6267 9643 6273
rect 9766 6264 9772 6276
rect 9824 6264 9830 6316
rect 14384 6313 14412 6344
rect 15286 6332 15292 6344
rect 15344 6332 15350 6384
rect 16546 6344 16580 6384
rect 16574 6332 16580 6344
rect 16632 6372 16638 6384
rect 16942 6372 16948 6384
rect 16632 6344 16948 6372
rect 16632 6332 16638 6344
rect 16942 6332 16948 6344
rect 17000 6332 17006 6384
rect 14369 6307 14427 6313
rect 14369 6273 14381 6307
rect 14415 6273 14427 6307
rect 14369 6267 14427 6273
rect 14550 6264 14556 6316
rect 14608 6264 14614 6316
rect 14642 6264 14648 6316
rect 14700 6304 14706 6316
rect 14829 6307 14887 6313
rect 14829 6304 14841 6307
rect 14700 6276 14841 6304
rect 14700 6264 14706 6276
rect 14829 6273 14841 6276
rect 14875 6273 14887 6307
rect 14829 6267 14887 6273
rect 16853 6307 16911 6313
rect 16853 6273 16865 6307
rect 16899 6304 16911 6307
rect 17218 6304 17224 6316
rect 16899 6276 17224 6304
rect 16899 6273 16911 6276
rect 16853 6267 16911 6273
rect 17218 6264 17224 6276
rect 17276 6264 17282 6316
rect 17862 6264 17868 6316
rect 17920 6304 17926 6316
rect 17956 6307 18014 6313
rect 17956 6304 17968 6307
rect 17920 6276 17968 6304
rect 17920 6264 17926 6276
rect 17956 6273 17968 6276
rect 18002 6273 18014 6307
rect 17956 6267 18014 6273
rect 18049 6307 18107 6313
rect 18049 6273 18061 6307
rect 18095 6304 18107 6307
rect 18598 6304 18604 6316
rect 18095 6276 18604 6304
rect 18095 6273 18107 6276
rect 18049 6267 18107 6273
rect 18598 6264 18604 6276
rect 18656 6264 18662 6316
rect 18782 6264 18788 6316
rect 18840 6264 18846 6316
rect 3418 6236 3424 6248
rect 3344 6208 3424 6236
rect 1670 6128 1676 6180
rect 1728 6168 1734 6180
rect 2222 6168 2228 6180
rect 1728 6140 2228 6168
rect 1728 6128 1734 6140
rect 2222 6128 2228 6140
rect 2280 6128 2286 6180
rect 3344 6177 3372 6208
rect 3418 6196 3424 6208
rect 3476 6196 3482 6248
rect 6914 6196 6920 6248
rect 6972 6236 6978 6248
rect 7558 6236 7564 6248
rect 6972 6208 7564 6236
rect 6972 6196 6978 6208
rect 7558 6196 7564 6208
rect 7616 6196 7622 6248
rect 7837 6239 7895 6245
rect 7837 6205 7849 6239
rect 7883 6236 7895 6239
rect 8846 6236 8852 6248
rect 7883 6208 8852 6236
rect 7883 6205 7895 6208
rect 7837 6199 7895 6205
rect 8846 6196 8852 6208
rect 8904 6196 8910 6248
rect 15010 6196 15016 6248
rect 15068 6196 15074 6248
rect 3329 6171 3387 6177
rect 3329 6137 3341 6171
rect 3375 6137 3387 6171
rect 3329 6131 3387 6137
rect 17494 6128 17500 6180
rect 17552 6168 17558 6180
rect 17681 6171 17739 6177
rect 17681 6168 17693 6171
rect 17552 6140 17693 6168
rect 17552 6128 17558 6140
rect 17681 6137 17693 6140
rect 17727 6137 17739 6171
rect 17681 6131 17739 6137
rect 1946 6060 1952 6112
rect 2004 6060 2010 6112
rect 13722 6060 13728 6112
rect 13780 6100 13786 6112
rect 13817 6103 13875 6109
rect 13817 6100 13829 6103
rect 13780 6072 13829 6100
rect 13780 6060 13786 6072
rect 13817 6069 13829 6072
rect 13863 6069 13875 6103
rect 13817 6063 13875 6069
rect 15473 6103 15531 6109
rect 15473 6069 15485 6103
rect 15519 6100 15531 6103
rect 17310 6100 17316 6112
rect 15519 6072 17316 6100
rect 15519 6069 15531 6072
rect 15473 6063 15531 6069
rect 17310 6060 17316 6072
rect 17368 6060 17374 6112
rect 1104 6010 19136 6032
rect 1104 5958 2350 6010
rect 2402 5958 2414 6010
rect 2466 5958 2478 6010
rect 2530 5958 2542 6010
rect 2594 5958 2606 6010
rect 2658 5958 19136 6010
rect 1104 5936 19136 5958
rect 2314 5856 2320 5908
rect 2372 5896 2378 5908
rect 3970 5896 3976 5908
rect 2372 5868 3976 5896
rect 2372 5856 2378 5868
rect 3970 5856 3976 5868
rect 4028 5856 4034 5908
rect 8294 5856 8300 5908
rect 8352 5896 8358 5908
rect 8389 5899 8447 5905
rect 8389 5896 8401 5899
rect 8352 5868 8401 5896
rect 8352 5856 8358 5868
rect 8389 5865 8401 5868
rect 8435 5865 8447 5899
rect 8389 5859 8447 5865
rect 8846 5856 8852 5908
rect 8904 5896 8910 5908
rect 8941 5899 8999 5905
rect 8941 5896 8953 5899
rect 8904 5868 8953 5896
rect 8904 5856 8910 5868
rect 8941 5865 8953 5868
rect 8987 5865 8999 5899
rect 8941 5859 8999 5865
rect 14550 5856 14556 5908
rect 14608 5896 14614 5908
rect 15577 5899 15635 5905
rect 15577 5896 15589 5899
rect 14608 5868 15589 5896
rect 14608 5856 14614 5868
rect 15577 5865 15589 5868
rect 15623 5896 15635 5899
rect 16393 5899 16451 5905
rect 16393 5896 16405 5899
rect 15623 5868 16405 5896
rect 15623 5865 15635 5868
rect 15577 5859 15635 5865
rect 16393 5865 16405 5868
rect 16439 5865 16451 5899
rect 16393 5859 16451 5865
rect 2225 5831 2283 5837
rect 2225 5797 2237 5831
rect 2271 5828 2283 5831
rect 2774 5828 2780 5840
rect 2271 5800 2780 5828
rect 2271 5797 2283 5800
rect 2225 5791 2283 5797
rect 2774 5788 2780 5800
rect 2832 5788 2838 5840
rect 3694 5788 3700 5840
rect 3752 5828 3758 5840
rect 3752 5800 4200 5828
rect 3752 5788 3758 5800
rect 1394 5720 1400 5772
rect 1452 5760 1458 5772
rect 2682 5760 2688 5772
rect 1452 5732 2688 5760
rect 1452 5720 1458 5732
rect 2682 5720 2688 5732
rect 2740 5760 2746 5772
rect 4065 5763 4123 5769
rect 4065 5760 4077 5763
rect 2740 5732 4077 5760
rect 2740 5720 2746 5732
rect 4065 5729 4077 5732
rect 4111 5729 4123 5763
rect 4172 5760 4200 5800
rect 8018 5788 8024 5840
rect 8076 5828 8082 5840
rect 8205 5831 8263 5837
rect 8205 5828 8217 5831
rect 8076 5800 8217 5828
rect 8076 5788 8082 5800
rect 8205 5797 8217 5800
rect 8251 5828 8263 5831
rect 8251 5800 9168 5828
rect 8251 5797 8263 5800
rect 8205 5791 8263 5797
rect 6822 5760 6828 5772
rect 4172 5732 6828 5760
rect 4065 5723 4123 5729
rect 6822 5720 6828 5732
rect 6880 5760 6886 5772
rect 6880 5732 8800 5760
rect 6880 5720 6886 5732
rect 8772 5704 8800 5732
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5692 1639 5695
rect 1857 5695 1915 5701
rect 1627 5664 1716 5692
rect 1627 5661 1639 5664
rect 1581 5655 1639 5661
rect 1397 5559 1455 5565
rect 1397 5525 1409 5559
rect 1443 5556 1455 5559
rect 1486 5556 1492 5568
rect 1443 5528 1492 5556
rect 1443 5525 1455 5528
rect 1397 5519 1455 5525
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 1688 5565 1716 5664
rect 1857 5661 1869 5695
rect 1903 5692 1915 5695
rect 2133 5695 2191 5701
rect 1903 5664 2084 5692
rect 1903 5661 1915 5664
rect 1857 5655 1915 5661
rect 1673 5559 1731 5565
rect 1673 5525 1685 5559
rect 1719 5525 1731 5559
rect 1673 5519 1731 5525
rect 1762 5516 1768 5568
rect 1820 5556 1826 5568
rect 1949 5559 2007 5565
rect 1949 5556 1961 5559
rect 1820 5528 1961 5556
rect 1820 5516 1826 5528
rect 1949 5525 1961 5528
rect 1995 5525 2007 5559
rect 2056 5556 2084 5664
rect 2133 5661 2145 5695
rect 2179 5692 2191 5695
rect 2222 5692 2228 5704
rect 2179 5664 2228 5692
rect 2179 5661 2191 5664
rect 2133 5655 2191 5661
rect 2222 5652 2228 5664
rect 2280 5652 2286 5704
rect 2314 5652 2320 5704
rect 2372 5652 2378 5704
rect 2409 5695 2467 5701
rect 2409 5661 2421 5695
rect 2455 5661 2467 5695
rect 2409 5655 2467 5661
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5692 2651 5695
rect 3510 5692 3516 5704
rect 2639 5664 3516 5692
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 2424 5624 2452 5655
rect 3510 5652 3516 5664
rect 3568 5652 3574 5704
rect 3786 5652 3792 5704
rect 3844 5652 3850 5704
rect 3970 5652 3976 5704
rect 4028 5652 4034 5704
rect 5902 5652 5908 5704
rect 5960 5692 5966 5704
rect 6089 5695 6147 5701
rect 6089 5692 6101 5695
rect 5960 5664 6101 5692
rect 5960 5652 5966 5664
rect 6089 5661 6101 5664
rect 6135 5692 6147 5695
rect 7006 5692 7012 5704
rect 6135 5664 7012 5692
rect 6135 5661 6147 5664
rect 6089 5655 6147 5661
rect 7006 5652 7012 5664
rect 7064 5652 7070 5704
rect 8110 5652 8116 5704
rect 8168 5652 8174 5704
rect 8754 5652 8760 5704
rect 8812 5652 8818 5704
rect 9140 5701 9168 5800
rect 10962 5788 10968 5840
rect 11020 5828 11026 5840
rect 11020 5800 12572 5828
rect 11020 5788 11026 5800
rect 9214 5720 9220 5772
rect 9272 5760 9278 5772
rect 11882 5760 11888 5772
rect 9272 5732 11888 5760
rect 9272 5720 9278 5732
rect 11882 5720 11888 5732
rect 11940 5760 11946 5772
rect 11940 5732 12480 5760
rect 11940 5720 11946 5732
rect 9125 5695 9183 5701
rect 9125 5661 9137 5695
rect 9171 5661 9183 5695
rect 9125 5655 9183 5661
rect 9306 5652 9312 5704
rect 9364 5652 9370 5704
rect 9401 5695 9459 5701
rect 9401 5661 9413 5695
rect 9447 5692 9459 5695
rect 9582 5692 9588 5704
rect 9447 5664 9588 5692
rect 9447 5661 9459 5664
rect 9401 5655 9459 5661
rect 9582 5652 9588 5664
rect 9640 5652 9646 5704
rect 9766 5652 9772 5704
rect 9824 5692 9830 5704
rect 10962 5692 10968 5704
rect 9824 5664 10968 5692
rect 9824 5652 9830 5664
rect 10962 5652 10968 5664
rect 11020 5692 11026 5704
rect 12452 5701 12480 5732
rect 12544 5701 12572 5800
rect 13722 5788 13728 5840
rect 13780 5788 13786 5840
rect 16022 5788 16028 5840
rect 16080 5788 16086 5840
rect 16408 5828 16436 5859
rect 16574 5856 16580 5908
rect 16632 5856 16638 5908
rect 18598 5856 18604 5908
rect 18656 5856 18662 5908
rect 16408 5800 16988 5828
rect 13740 5760 13768 5788
rect 15562 5760 15568 5772
rect 13740 5732 15568 5760
rect 15562 5720 15568 5732
rect 15620 5760 15626 5772
rect 15841 5763 15899 5769
rect 15841 5760 15853 5763
rect 15620 5732 15853 5760
rect 15620 5720 15626 5732
rect 15841 5729 15853 5732
rect 15887 5760 15899 5763
rect 16853 5763 16911 5769
rect 16853 5760 16865 5763
rect 15887 5732 16865 5760
rect 15887 5729 15899 5732
rect 15841 5723 15899 5729
rect 16853 5729 16865 5732
rect 16899 5729 16911 5763
rect 16960 5760 16988 5800
rect 17862 5760 17868 5772
rect 16960 5732 17868 5760
rect 16853 5723 16911 5729
rect 17862 5720 17868 5732
rect 17920 5720 17926 5772
rect 11057 5695 11115 5701
rect 11057 5692 11069 5695
rect 11020 5664 11069 5692
rect 11020 5652 11026 5664
rect 11057 5661 11069 5664
rect 11103 5661 11115 5695
rect 11057 5655 11115 5661
rect 12344 5695 12402 5701
rect 12344 5661 12356 5695
rect 12390 5661 12402 5695
rect 12344 5655 12402 5661
rect 12437 5695 12495 5701
rect 12437 5661 12449 5695
rect 12483 5661 12495 5695
rect 12437 5655 12495 5661
rect 12529 5695 12587 5701
rect 12529 5661 12541 5695
rect 12575 5692 12587 5695
rect 13446 5692 13452 5704
rect 12575 5664 13452 5692
rect 12575 5661 12587 5664
rect 12529 5655 12587 5661
rect 3602 5624 3608 5636
rect 2424 5596 3608 5624
rect 3602 5584 3608 5596
rect 3660 5584 3666 5636
rect 3881 5627 3939 5633
rect 3881 5593 3893 5627
rect 3927 5624 3939 5627
rect 4341 5627 4399 5633
rect 4341 5624 4353 5627
rect 3927 5596 4353 5624
rect 3927 5593 3939 5596
rect 3881 5587 3939 5593
rect 4341 5593 4353 5596
rect 4387 5593 4399 5627
rect 5997 5627 6055 5633
rect 5997 5624 6009 5627
rect 5566 5596 6009 5624
rect 4341 5587 4399 5593
rect 5997 5593 6009 5596
rect 6043 5593 6055 5627
rect 12360 5624 12388 5655
rect 13446 5652 13452 5664
rect 13504 5692 13510 5704
rect 13725 5695 13783 5701
rect 13725 5692 13737 5695
rect 13504 5664 13737 5692
rect 13504 5652 13510 5664
rect 13725 5661 13737 5664
rect 13771 5692 13783 5695
rect 14274 5692 14280 5704
rect 13771 5664 14280 5692
rect 13771 5661 13783 5664
rect 13725 5655 13783 5661
rect 14274 5652 14280 5664
rect 14332 5652 14338 5704
rect 13262 5624 13268 5636
rect 12360 5596 13268 5624
rect 5997 5587 6055 5593
rect 13262 5584 13268 5596
rect 13320 5584 13326 5636
rect 13817 5627 13875 5633
rect 13817 5593 13829 5627
rect 13863 5624 13875 5627
rect 13863 5596 14398 5624
rect 13863 5593 13875 5596
rect 13817 5587 13875 5593
rect 17126 5584 17132 5636
rect 17184 5584 17190 5636
rect 18138 5584 18144 5636
rect 18196 5584 18202 5636
rect 2774 5556 2780 5568
rect 2056 5528 2780 5556
rect 1949 5519 2007 5525
rect 2774 5516 2780 5528
rect 2832 5516 2838 5568
rect 5810 5516 5816 5568
rect 5868 5516 5874 5568
rect 6825 5559 6883 5565
rect 6825 5525 6837 5559
rect 6871 5556 6883 5559
rect 6914 5556 6920 5568
rect 6871 5528 6920 5556
rect 6871 5525 6883 5528
rect 6825 5519 6883 5525
rect 6914 5516 6920 5528
rect 6972 5516 6978 5568
rect 8389 5559 8447 5565
rect 8389 5525 8401 5559
rect 8435 5556 8447 5559
rect 8570 5556 8576 5568
rect 8435 5528 8576 5556
rect 8435 5525 8447 5528
rect 8389 5519 8447 5525
rect 8570 5516 8576 5528
rect 8628 5516 8634 5568
rect 10962 5516 10968 5568
rect 11020 5516 11026 5568
rect 12066 5516 12072 5568
rect 12124 5516 12130 5568
rect 12526 5516 12532 5568
rect 12584 5556 12590 5568
rect 12621 5559 12679 5565
rect 12621 5556 12633 5559
rect 12584 5528 12633 5556
rect 12584 5516 12590 5528
rect 12621 5525 12633 5528
rect 12667 5525 12679 5559
rect 12621 5519 12679 5525
rect 14093 5559 14151 5565
rect 14093 5525 14105 5559
rect 14139 5556 14151 5559
rect 14734 5556 14740 5568
rect 14139 5528 14740 5556
rect 14139 5525 14151 5528
rect 14093 5519 14151 5525
rect 14734 5516 14740 5528
rect 14792 5516 14798 5568
rect 16393 5559 16451 5565
rect 16393 5525 16405 5559
rect 16439 5556 16451 5559
rect 16482 5556 16488 5568
rect 16439 5528 16488 5556
rect 16439 5525 16451 5528
rect 16393 5519 16451 5525
rect 16482 5516 16488 5528
rect 16540 5516 16546 5568
rect 1104 5466 19136 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 19136 5466
rect 1104 5392 19136 5414
rect 2774 5312 2780 5364
rect 2832 5352 2838 5364
rect 3237 5355 3295 5361
rect 3237 5352 3249 5355
rect 2832 5324 3249 5352
rect 2832 5312 2838 5324
rect 3237 5321 3249 5324
rect 3283 5321 3295 5355
rect 3237 5315 3295 5321
rect 3510 5312 3516 5364
rect 3568 5312 3574 5364
rect 5810 5352 5816 5364
rect 5092 5324 5816 5352
rect 1762 5244 1768 5296
rect 1820 5244 1826 5296
rect 3970 5284 3976 5296
rect 3620 5256 3976 5284
rect 3620 5228 3648 5256
rect 3970 5244 3976 5256
rect 4028 5244 4034 5296
rect 1394 5176 1400 5228
rect 1452 5216 1458 5228
rect 1489 5219 1547 5225
rect 1489 5216 1501 5219
rect 1452 5188 1501 5216
rect 1452 5176 1458 5188
rect 1489 5185 1501 5188
rect 1535 5185 1547 5219
rect 1489 5179 1547 5185
rect 2866 5176 2872 5228
rect 2924 5176 2930 5228
rect 3602 5176 3608 5228
rect 3660 5176 3666 5228
rect 3786 5176 3792 5228
rect 3844 5176 3850 5228
rect 4801 5219 4859 5225
rect 4801 5185 4813 5219
rect 4847 5185 4859 5219
rect 4801 5179 4859 5185
rect 4955 5219 5013 5225
rect 4955 5185 4967 5219
rect 5001 5216 5013 5219
rect 5092 5216 5120 5324
rect 5810 5312 5816 5324
rect 5868 5312 5874 5364
rect 9030 5352 9036 5364
rect 7300 5324 9036 5352
rect 5169 5287 5227 5293
rect 5169 5253 5181 5287
rect 5215 5284 5227 5287
rect 5445 5287 5503 5293
rect 5445 5284 5457 5287
rect 5215 5256 5457 5284
rect 5215 5253 5227 5256
rect 5169 5247 5227 5253
rect 5445 5253 5457 5256
rect 5491 5253 5503 5287
rect 5445 5247 5503 5253
rect 5994 5244 6000 5296
rect 6052 5244 6058 5296
rect 7300 5284 7328 5324
rect 9030 5312 9036 5324
rect 9088 5312 9094 5364
rect 9493 5355 9551 5361
rect 9493 5321 9505 5355
rect 9539 5352 9551 5355
rect 11238 5352 11244 5364
rect 9539 5324 11244 5352
rect 9539 5321 9551 5324
rect 9493 5315 9551 5321
rect 11238 5312 11244 5324
rect 11296 5312 11302 5364
rect 13262 5312 13268 5364
rect 13320 5312 13326 5364
rect 15010 5312 15016 5364
rect 15068 5312 15074 5364
rect 17037 5355 17095 5361
rect 17037 5321 17049 5355
rect 17083 5352 17095 5355
rect 17126 5352 17132 5364
rect 17083 5324 17132 5352
rect 17083 5321 17095 5324
rect 17037 5315 17095 5321
rect 17126 5312 17132 5324
rect 17184 5312 17190 5364
rect 17957 5355 18015 5361
rect 17957 5321 17969 5355
rect 18003 5352 18015 5355
rect 18138 5352 18144 5364
rect 18003 5324 18144 5352
rect 18003 5321 18015 5324
rect 17957 5315 18015 5321
rect 18138 5312 18144 5324
rect 18196 5312 18202 5364
rect 18782 5312 18788 5364
rect 18840 5312 18846 5364
rect 6840 5256 7328 5284
rect 5001 5188 5120 5216
rect 5001 5185 5013 5188
rect 4955 5179 5013 5185
rect 2222 5108 2228 5160
rect 2280 5148 2286 5160
rect 3804 5148 3832 5176
rect 2280 5120 3832 5148
rect 2280 5108 2286 5120
rect 3329 5083 3387 5089
rect 3329 5049 3341 5083
rect 3375 5080 3387 5083
rect 4062 5080 4068 5092
rect 3375 5052 4068 5080
rect 3375 5049 3387 5052
rect 3329 5043 3387 5049
rect 4062 5040 4068 5052
rect 4120 5040 4126 5092
rect 4816 5012 4844 5179
rect 5350 5108 5356 5160
rect 5408 5108 5414 5160
rect 6840 5012 6868 5256
rect 7006 5176 7012 5228
rect 7064 5176 7070 5228
rect 7300 5225 7328 5256
rect 8018 5244 8024 5296
rect 8076 5244 8082 5296
rect 9582 5284 9588 5296
rect 9246 5256 9588 5284
rect 9582 5244 9588 5256
rect 9640 5244 9646 5296
rect 10962 5284 10968 5296
rect 10626 5256 10968 5284
rect 10962 5244 10968 5256
rect 11020 5244 11026 5296
rect 11422 5244 11428 5296
rect 11480 5284 11486 5296
rect 11793 5287 11851 5293
rect 11793 5284 11805 5287
rect 11480 5256 11805 5284
rect 11480 5244 11486 5256
rect 11793 5253 11805 5256
rect 11839 5253 11851 5287
rect 11793 5247 11851 5253
rect 12526 5244 12532 5296
rect 12584 5244 12590 5296
rect 14274 5244 14280 5296
rect 14332 5284 14338 5296
rect 14332 5256 15424 5284
rect 14332 5244 14338 5256
rect 7285 5219 7343 5225
rect 7285 5185 7297 5219
rect 7331 5185 7343 5219
rect 7285 5179 7343 5185
rect 7439 5219 7497 5225
rect 7439 5185 7451 5219
rect 7485 5216 7497 5219
rect 7650 5216 7656 5228
rect 7485 5188 7656 5216
rect 7485 5185 7497 5188
rect 7439 5179 7497 5185
rect 7650 5176 7656 5188
rect 7708 5176 7714 5228
rect 14645 5219 14703 5225
rect 14645 5185 14657 5219
rect 14691 5185 14703 5219
rect 14645 5179 14703 5185
rect 6914 5108 6920 5160
rect 6972 5148 6978 5160
rect 7745 5151 7803 5157
rect 7745 5148 7757 5151
rect 6972 5120 7757 5148
rect 6972 5108 6978 5120
rect 7745 5117 7757 5120
rect 7791 5117 7803 5151
rect 7745 5111 7803 5117
rect 11054 5108 11060 5160
rect 11112 5108 11118 5160
rect 11333 5151 11391 5157
rect 11333 5117 11345 5151
rect 11379 5148 11391 5151
rect 11514 5148 11520 5160
rect 11379 5120 11520 5148
rect 11379 5117 11391 5120
rect 11333 5111 11391 5117
rect 11514 5108 11520 5120
rect 11572 5108 11578 5160
rect 14660 5148 14688 5179
rect 14734 5176 14740 5228
rect 14792 5216 14798 5228
rect 15396 5225 15424 5256
rect 17218 5244 17224 5296
rect 17276 5284 17282 5296
rect 17276 5256 17908 5284
rect 17276 5244 17282 5256
rect 15381 5219 15439 5225
rect 14792 5188 14837 5216
rect 14792 5176 14798 5188
rect 15381 5185 15393 5219
rect 15427 5216 15439 5219
rect 15427 5188 16574 5216
rect 15427 5185 15439 5188
rect 15381 5179 15439 5185
rect 15930 5148 15936 5160
rect 14660 5120 15936 5148
rect 15930 5108 15936 5120
rect 15988 5108 15994 5160
rect 16546 5148 16574 5188
rect 17126 5176 17132 5228
rect 17184 5216 17190 5228
rect 17313 5219 17371 5225
rect 17313 5216 17325 5219
rect 17184 5188 17325 5216
rect 17184 5176 17190 5188
rect 17313 5185 17325 5188
rect 17359 5185 17371 5219
rect 17313 5179 17371 5185
rect 17405 5219 17463 5225
rect 17405 5185 17417 5219
rect 17451 5185 17463 5219
rect 17405 5179 17463 5185
rect 17218 5148 17224 5160
rect 16546 5120 17224 5148
rect 17218 5108 17224 5120
rect 17276 5108 17282 5160
rect 17310 5040 17316 5092
rect 17368 5080 17374 5092
rect 17420 5080 17448 5179
rect 17494 5176 17500 5228
rect 17552 5176 17558 5228
rect 17678 5176 17684 5228
rect 17736 5176 17742 5228
rect 17880 5225 17908 5256
rect 17865 5219 17923 5225
rect 17865 5185 17877 5219
rect 17911 5185 17923 5219
rect 17865 5179 17923 5185
rect 18506 5176 18512 5228
rect 18564 5216 18570 5228
rect 18601 5219 18659 5225
rect 18601 5216 18613 5219
rect 18564 5188 18613 5216
rect 18564 5176 18570 5188
rect 18601 5185 18613 5188
rect 18647 5185 18659 5219
rect 18601 5179 18659 5185
rect 18138 5080 18144 5092
rect 17368 5052 18144 5080
rect 17368 5040 17374 5052
rect 18138 5040 18144 5052
rect 18196 5040 18202 5092
rect 4816 4984 6868 5012
rect 7006 4972 7012 5024
rect 7064 5012 7070 5024
rect 7101 5015 7159 5021
rect 7101 5012 7113 5015
rect 7064 4984 7113 5012
rect 7064 4972 7070 4984
rect 7101 4981 7113 4984
rect 7147 4981 7159 5015
rect 7101 4975 7159 4981
rect 7466 4972 7472 5024
rect 7524 4972 7530 5024
rect 9585 5015 9643 5021
rect 9585 4981 9597 5015
rect 9631 5012 9643 5015
rect 10686 5012 10692 5024
rect 9631 4984 10692 5012
rect 9631 4981 9643 4984
rect 9585 4975 9643 4981
rect 10686 4972 10692 4984
rect 10744 4972 10750 5024
rect 15378 4972 15384 5024
rect 15436 5012 15442 5024
rect 15473 5015 15531 5021
rect 15473 5012 15485 5015
rect 15436 4984 15485 5012
rect 15436 4972 15442 4984
rect 15473 4981 15485 4984
rect 15519 4981 15531 5015
rect 15473 4975 15531 4981
rect 17126 4972 17132 5024
rect 17184 5012 17190 5024
rect 17862 5012 17868 5024
rect 17184 4984 17868 5012
rect 17184 4972 17190 4984
rect 17862 4972 17868 4984
rect 17920 5012 17926 5024
rect 18046 5012 18052 5024
rect 17920 4984 18052 5012
rect 17920 4972 17926 4984
rect 18046 4972 18052 4984
rect 18104 4972 18110 5024
rect 1104 4922 19136 4944
rect 1104 4870 2350 4922
rect 2402 4870 2414 4922
rect 2466 4870 2478 4922
rect 2530 4870 2542 4922
rect 2594 4870 2606 4922
rect 2658 4870 19136 4922
rect 1104 4848 19136 4870
rect 2593 4811 2651 4817
rect 2593 4777 2605 4811
rect 2639 4808 2651 4811
rect 2866 4808 2872 4820
rect 2639 4780 2872 4808
rect 2639 4777 2651 4780
rect 2593 4771 2651 4777
rect 2866 4768 2872 4780
rect 2924 4768 2930 4820
rect 3786 4768 3792 4820
rect 3844 4808 3850 4820
rect 3927 4811 3985 4817
rect 3927 4808 3939 4811
rect 3844 4780 3939 4808
rect 3844 4768 3850 4780
rect 3927 4777 3939 4780
rect 3973 4777 3985 4811
rect 3927 4771 3985 4777
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 7745 4811 7803 4817
rect 7745 4808 7757 4811
rect 7708 4780 7757 4808
rect 7708 4768 7714 4780
rect 7745 4777 7757 4780
rect 7791 4777 7803 4811
rect 7745 4771 7803 4777
rect 9582 4768 9588 4820
rect 9640 4768 9646 4820
rect 11054 4768 11060 4820
rect 11112 4808 11118 4820
rect 11149 4811 11207 4817
rect 11149 4808 11161 4811
rect 11112 4780 11161 4808
rect 11112 4768 11118 4780
rect 11149 4777 11161 4780
rect 11195 4777 11207 4811
rect 11149 4771 11207 4777
rect 16390 4768 16396 4820
rect 16448 4768 16454 4820
rect 1946 4632 1952 4684
rect 2004 4672 2010 4684
rect 2869 4675 2927 4681
rect 2004 4644 2820 4672
rect 2004 4632 2010 4644
rect 842 4564 848 4616
rect 900 4604 906 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 900 4576 1409 4604
rect 900 4564 906 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 2130 4564 2136 4616
rect 2188 4604 2194 4616
rect 2792 4613 2820 4644
rect 2869 4641 2881 4675
rect 2915 4672 2927 4675
rect 3602 4672 3608 4684
rect 2915 4644 3608 4672
rect 2915 4641 2927 4644
rect 2869 4635 2927 4641
rect 3602 4632 3608 4644
rect 3660 4672 3666 4684
rect 4065 4675 4123 4681
rect 4065 4672 4077 4675
rect 3660 4644 4077 4672
rect 3660 4632 3666 4644
rect 4065 4641 4077 4644
rect 4111 4641 4123 4675
rect 6914 4672 6920 4684
rect 4065 4635 4123 4641
rect 6012 4644 6920 4672
rect 2501 4607 2559 4613
rect 2501 4604 2513 4607
rect 2188 4576 2513 4604
rect 2188 4564 2194 4576
rect 2501 4573 2513 4576
rect 2547 4573 2559 4607
rect 2501 4567 2559 4573
rect 2777 4607 2835 4613
rect 2777 4573 2789 4607
rect 2823 4573 2835 4607
rect 2777 4567 2835 4573
rect 3694 4564 3700 4616
rect 3752 4604 3758 4616
rect 3789 4607 3847 4613
rect 3789 4604 3801 4607
rect 3752 4576 3801 4604
rect 3752 4564 3758 4576
rect 3789 4573 3801 4576
rect 3835 4573 3847 4607
rect 3789 4567 3847 4573
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4604 4307 4607
rect 5350 4604 5356 4616
rect 4295 4576 5356 4604
rect 4295 4573 4307 4576
rect 4249 4567 4307 4573
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 5534 4564 5540 4616
rect 5592 4604 5598 4616
rect 6012 4613 6040 4644
rect 6914 4632 6920 4644
rect 6972 4632 6978 4684
rect 11977 4675 12035 4681
rect 11977 4672 11989 4675
rect 10704 4644 11989 4672
rect 10704 4616 10732 4644
rect 11977 4641 11989 4644
rect 12023 4641 12035 4675
rect 11977 4635 12035 4641
rect 12066 4632 12072 4684
rect 12124 4672 12130 4684
rect 12161 4675 12219 4681
rect 12161 4672 12173 4675
rect 12124 4644 12173 4672
rect 12124 4632 12130 4644
rect 12161 4641 12173 4644
rect 12207 4641 12219 4675
rect 12161 4635 12219 4641
rect 16117 4675 16175 4681
rect 16117 4641 16129 4675
rect 16163 4672 16175 4675
rect 16163 4644 16344 4672
rect 16163 4641 16175 4644
rect 16117 4635 16175 4641
rect 5997 4607 6055 4613
rect 5997 4604 6009 4607
rect 5592 4576 6009 4604
rect 5592 4564 5598 4576
rect 5997 4573 6009 4576
rect 6043 4573 6055 4607
rect 5997 4567 6055 4573
rect 9677 4607 9735 4613
rect 9677 4573 9689 4607
rect 9723 4604 9735 4607
rect 9766 4604 9772 4616
rect 9723 4576 9772 4604
rect 9723 4573 9735 4576
rect 9677 4567 9735 4573
rect 9766 4564 9772 4576
rect 9824 4564 9830 4616
rect 10686 4564 10692 4616
rect 10744 4564 10750 4616
rect 10965 4607 11023 4613
rect 10965 4573 10977 4607
rect 11011 4604 11023 4607
rect 11146 4604 11152 4616
rect 11011 4576 11152 4604
rect 11011 4573 11023 4576
rect 10965 4567 11023 4573
rect 11146 4564 11152 4576
rect 11204 4564 11210 4616
rect 11241 4607 11299 4613
rect 11241 4573 11253 4607
rect 11287 4573 11299 4607
rect 11241 4567 11299 4573
rect 2038 4496 2044 4548
rect 2096 4536 2102 4548
rect 2225 4539 2283 4545
rect 2225 4536 2237 4539
rect 2096 4508 2237 4536
rect 2096 4496 2102 4508
rect 2225 4505 2237 4508
rect 2271 4536 2283 4539
rect 3712 4536 3740 4564
rect 2271 4508 3740 4536
rect 6273 4539 6331 4545
rect 2271 4505 2283 4508
rect 2225 4499 2283 4505
rect 6273 4505 6285 4539
rect 6319 4505 6331 4539
rect 6273 4499 6331 4505
rect 4154 4428 4160 4480
rect 4212 4428 4218 4480
rect 6288 4468 6316 4499
rect 7006 4496 7012 4548
rect 7064 4496 7070 4548
rect 8662 4496 8668 4548
rect 8720 4536 8726 4548
rect 11256 4536 11284 4567
rect 11422 4564 11428 4616
rect 11480 4564 11486 4616
rect 13722 4564 13728 4616
rect 13780 4604 13786 4616
rect 14369 4607 14427 4613
rect 14369 4604 14381 4607
rect 13780 4576 14381 4604
rect 13780 4564 13786 4576
rect 14369 4573 14381 4576
rect 14415 4573 14427 4607
rect 14369 4567 14427 4573
rect 15930 4564 15936 4616
rect 15988 4604 15994 4616
rect 16316 4613 16344 4644
rect 16209 4607 16267 4613
rect 16209 4604 16221 4607
rect 15988 4576 16221 4604
rect 15988 4564 15994 4576
rect 16209 4573 16221 4576
rect 16255 4573 16267 4607
rect 16209 4567 16267 4573
rect 16302 4607 16360 4613
rect 16302 4573 16314 4607
rect 16348 4573 16360 4607
rect 16302 4567 16360 4573
rect 17770 4564 17776 4616
rect 17828 4604 17834 4616
rect 18079 4607 18137 4613
rect 18079 4604 18091 4607
rect 17828 4576 18091 4604
rect 17828 4564 17834 4576
rect 18079 4573 18091 4576
rect 18125 4573 18137 4607
rect 18079 4567 18137 4573
rect 18230 4564 18236 4616
rect 18288 4564 18294 4616
rect 18322 4564 18328 4616
rect 18380 4604 18386 4616
rect 18601 4607 18659 4613
rect 18601 4604 18613 4607
rect 18380 4576 18613 4604
rect 18380 4564 18386 4576
rect 18601 4573 18613 4576
rect 18647 4573 18659 4607
rect 18601 4567 18659 4573
rect 11330 4536 11336 4548
rect 8720 4508 11336 4536
rect 8720 4496 8726 4508
rect 11330 4496 11336 4508
rect 11388 4496 11394 4548
rect 14645 4539 14703 4545
rect 14645 4505 14657 4539
rect 14691 4505 14703 4539
rect 14645 4499 14703 4505
rect 6638 4468 6644 4480
rect 6288 4440 6644 4468
rect 6638 4428 6644 4440
rect 6696 4428 6702 4480
rect 10781 4471 10839 4477
rect 10781 4437 10793 4471
rect 10827 4468 10839 4471
rect 11241 4471 11299 4477
rect 11241 4468 11253 4471
rect 10827 4440 11253 4468
rect 10827 4437 10839 4440
rect 10781 4431 10839 4437
rect 11241 4437 11253 4440
rect 11287 4437 11299 4471
rect 11241 4431 11299 4437
rect 12618 4428 12624 4480
rect 12676 4428 12682 4480
rect 14660 4468 14688 4499
rect 15378 4496 15384 4548
rect 15436 4496 15442 4548
rect 16574 4468 16580 4480
rect 14660 4440 16580 4468
rect 16574 4428 16580 4440
rect 16632 4428 16638 4480
rect 17678 4428 17684 4480
rect 17736 4468 17742 4480
rect 17865 4471 17923 4477
rect 17865 4468 17877 4471
rect 17736 4440 17877 4468
rect 17736 4428 17742 4440
rect 17865 4437 17877 4440
rect 17911 4437 17923 4471
rect 17865 4431 17923 4437
rect 18782 4428 18788 4480
rect 18840 4428 18846 4480
rect 1104 4378 19136 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 19136 4378
rect 1104 4304 19136 4326
rect 4154 4224 4160 4276
rect 4212 4224 4218 4276
rect 5261 4267 5319 4273
rect 5261 4233 5273 4267
rect 5307 4264 5319 4267
rect 5350 4264 5356 4276
rect 5307 4236 5356 4264
rect 5307 4233 5319 4236
rect 5261 4227 5319 4233
rect 5350 4224 5356 4236
rect 5408 4224 5414 4276
rect 11330 4224 11336 4276
rect 11388 4264 11394 4276
rect 11388 4236 12848 4264
rect 11388 4224 11394 4236
rect 2222 4196 2228 4208
rect 2148 4168 2228 4196
rect 1670 4088 1676 4140
rect 1728 4088 1734 4140
rect 2038 4088 2044 4140
rect 2096 4088 2102 4140
rect 1581 4063 1639 4069
rect 1581 4029 1593 4063
rect 1627 4060 1639 4063
rect 1946 4060 1952 4072
rect 1627 4032 1952 4060
rect 1627 4029 1639 4032
rect 1581 4023 1639 4029
rect 1946 4020 1952 4032
rect 2004 4020 2010 4072
rect 2148 4060 2176 4168
rect 2222 4156 2228 4168
rect 2280 4156 2286 4208
rect 4172 4196 4200 4224
rect 8110 4196 8116 4208
rect 3528 4168 4200 4196
rect 6564 4168 8116 4196
rect 3234 4128 3240 4140
rect 2056 4032 2176 4060
rect 2240 4100 3240 4128
rect 2056 3933 2084 4032
rect 2240 4001 2268 4100
rect 3234 4088 3240 4100
rect 3292 4088 3298 4140
rect 3421 4131 3479 4137
rect 3421 4097 3433 4131
rect 3467 4128 3479 4131
rect 3528 4128 3556 4168
rect 5445 4131 5503 4137
rect 5445 4128 5457 4131
rect 3467 4100 3556 4128
rect 4922 4100 5457 4128
rect 3467 4097 3479 4100
rect 3421 4091 3479 4097
rect 5445 4097 5457 4100
rect 5491 4097 5503 4131
rect 5445 4091 5503 4097
rect 5537 4131 5595 4137
rect 5537 4097 5549 4131
rect 5583 4128 5595 4131
rect 5718 4128 5724 4140
rect 5583 4100 5724 4128
rect 5583 4097 5595 4100
rect 5537 4091 5595 4097
rect 5718 4088 5724 4100
rect 5776 4128 5782 4140
rect 6564 4128 6592 4168
rect 7116 4140 7144 4168
rect 8110 4156 8116 4168
rect 8168 4156 8174 4208
rect 12452 4168 12756 4196
rect 5776 4100 6592 4128
rect 5776 4088 5782 4100
rect 6638 4088 6644 4140
rect 6696 4088 6702 4140
rect 6822 4088 6828 4140
rect 6880 4088 6886 4140
rect 6917 4131 6975 4137
rect 6917 4097 6929 4131
rect 6963 4097 6975 4131
rect 6917 4091 6975 4097
rect 2682 4020 2688 4072
rect 2740 4060 2746 4072
rect 3513 4063 3571 4069
rect 3513 4060 3525 4063
rect 2740 4032 3525 4060
rect 2740 4020 2746 4032
rect 3513 4029 3525 4032
rect 3559 4029 3571 4063
rect 3789 4063 3847 4069
rect 3789 4060 3801 4063
rect 3513 4023 3571 4029
rect 3620 4032 3801 4060
rect 2225 3995 2283 4001
rect 2225 3961 2237 3995
rect 2271 3961 2283 3995
rect 2225 3955 2283 3961
rect 3329 3995 3387 4001
rect 3329 3961 3341 3995
rect 3375 3992 3387 3995
rect 3620 3992 3648 4032
rect 3789 4029 3801 4032
rect 3835 4029 3847 4063
rect 6932 4060 6960 4091
rect 7098 4088 7104 4140
rect 7156 4128 7162 4140
rect 7193 4131 7251 4137
rect 7193 4128 7205 4131
rect 7156 4100 7205 4128
rect 7156 4088 7162 4100
rect 7193 4097 7205 4100
rect 7239 4097 7251 4131
rect 7193 4091 7251 4097
rect 7466 4088 7472 4140
rect 7524 4128 7530 4140
rect 7745 4131 7803 4137
rect 7745 4128 7757 4131
rect 7524 4100 7757 4128
rect 7524 4088 7530 4100
rect 7745 4097 7757 4100
rect 7791 4097 7803 4131
rect 7745 4091 7803 4097
rect 8846 4088 8852 4140
rect 8904 4137 8910 4140
rect 8904 4131 8937 4137
rect 8925 4097 8937 4131
rect 8904 4091 8937 4097
rect 9033 4131 9091 4137
rect 9033 4097 9045 4131
rect 9079 4128 9091 4131
rect 10686 4128 10692 4140
rect 9079 4100 10692 4128
rect 9079 4097 9091 4100
rect 9033 4091 9091 4097
rect 8904 4088 8910 4091
rect 10686 4088 10692 4100
rect 10744 4088 10750 4140
rect 11882 4088 11888 4140
rect 11940 4128 11946 4140
rect 12452 4128 12480 4168
rect 11940 4100 12480 4128
rect 12529 4131 12587 4137
rect 11940 4088 11946 4100
rect 12529 4097 12541 4131
rect 12575 4097 12587 4131
rect 12529 4091 12587 4097
rect 7282 4060 7288 4072
rect 6932 4032 7288 4060
rect 3789 4023 3847 4029
rect 7282 4020 7288 4032
rect 7340 4060 7346 4072
rect 7561 4063 7619 4069
rect 7561 4060 7573 4063
rect 7340 4032 7573 4060
rect 7340 4020 7346 4032
rect 7561 4029 7573 4032
rect 7607 4029 7619 4063
rect 7561 4023 7619 4029
rect 11974 4020 11980 4072
rect 12032 4060 12038 4072
rect 12544 4060 12572 4091
rect 12618 4088 12624 4140
rect 12676 4088 12682 4140
rect 12728 4137 12756 4168
rect 12713 4131 12771 4137
rect 12713 4097 12725 4131
rect 12759 4097 12771 4131
rect 12820 4128 12848 4236
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 12820 4100 12909 4128
rect 12713 4091 12771 4097
rect 12897 4097 12909 4100
rect 12943 4128 12955 4131
rect 12986 4128 12992 4140
rect 12943 4100 12992 4128
rect 12943 4097 12955 4100
rect 12897 4091 12955 4097
rect 12986 4088 12992 4100
rect 13044 4088 13050 4140
rect 13446 4088 13452 4140
rect 13504 4088 13510 4140
rect 15194 4088 15200 4140
rect 15252 4088 15258 4140
rect 15381 4131 15439 4137
rect 15381 4097 15393 4131
rect 15427 4097 15439 4131
rect 15381 4091 15439 4097
rect 15473 4131 15531 4137
rect 15473 4097 15485 4131
rect 15519 4128 15531 4131
rect 16025 4131 16083 4137
rect 15519 4100 15884 4128
rect 15519 4097 15531 4100
rect 15473 4091 15531 4097
rect 12032 4032 12572 4060
rect 12636 4060 12664 4088
rect 12636 4032 12940 4060
rect 12032 4020 12038 4032
rect 12912 4004 12940 4032
rect 3375 3964 3648 3992
rect 3375 3961 3387 3964
rect 3329 3955 3387 3961
rect 8294 3952 8300 4004
rect 8352 3992 8358 4004
rect 8665 3995 8723 4001
rect 8665 3992 8677 3995
rect 8352 3964 8677 3992
rect 8352 3952 8358 3964
rect 8665 3961 8677 3964
rect 8711 3961 8723 3995
rect 8665 3955 8723 3961
rect 12894 3952 12900 4004
rect 12952 3952 12958 4004
rect 15396 3992 15424 4091
rect 15856 4072 15884 4100
rect 16025 4097 16037 4131
rect 16071 4128 16083 4131
rect 16390 4128 16396 4140
rect 16071 4100 16396 4128
rect 16071 4097 16083 4100
rect 16025 4091 16083 4097
rect 16390 4088 16396 4100
rect 16448 4088 16454 4140
rect 18414 4088 18420 4140
rect 18472 4088 18478 4140
rect 15838 4020 15844 4072
rect 15896 4020 15902 4072
rect 17034 4020 17040 4072
rect 17092 4020 17098 4072
rect 17310 4020 17316 4072
rect 17368 4020 17374 4072
rect 15930 3992 15936 4004
rect 15396 3964 15936 3992
rect 15930 3952 15936 3964
rect 15988 3952 15994 4004
rect 2041 3927 2099 3933
rect 2041 3893 2053 3927
rect 2087 3893 2099 3927
rect 2041 3887 2099 3893
rect 5810 3884 5816 3936
rect 5868 3924 5874 3936
rect 6457 3927 6515 3933
rect 6457 3924 6469 3927
rect 5868 3896 6469 3924
rect 5868 3884 5874 3896
rect 6457 3893 6469 3896
rect 6503 3893 6515 3927
rect 6457 3887 6515 3893
rect 7098 3884 7104 3936
rect 7156 3884 7162 3936
rect 8205 3927 8263 3933
rect 8205 3893 8217 3927
rect 8251 3924 8263 3927
rect 8386 3924 8392 3936
rect 8251 3896 8392 3924
rect 8251 3893 8263 3896
rect 8205 3887 8263 3893
rect 8386 3884 8392 3896
rect 8444 3884 8450 3936
rect 12250 3884 12256 3936
rect 12308 3884 12314 3936
rect 13357 3927 13415 3933
rect 13357 3893 13369 3927
rect 13403 3924 13415 3927
rect 13446 3924 13452 3936
rect 13403 3896 13452 3924
rect 13403 3893 13415 3896
rect 13357 3887 13415 3893
rect 13446 3884 13452 3896
rect 13504 3884 13510 3936
rect 14366 3884 14372 3936
rect 14424 3924 14430 3936
rect 15013 3927 15071 3933
rect 15013 3924 15025 3927
rect 14424 3896 15025 3924
rect 14424 3884 14430 3896
rect 15013 3893 15025 3896
rect 15059 3893 15071 3927
rect 15013 3887 15071 3893
rect 16485 3927 16543 3933
rect 16485 3893 16497 3927
rect 16531 3924 16543 3927
rect 17494 3924 17500 3936
rect 16531 3896 17500 3924
rect 16531 3893 16543 3896
rect 16485 3887 16543 3893
rect 17494 3884 17500 3896
rect 17552 3884 17558 3936
rect 18782 3884 18788 3936
rect 18840 3884 18846 3936
rect 1104 3834 19136 3856
rect 1104 3782 2350 3834
rect 2402 3782 2414 3834
rect 2466 3782 2478 3834
rect 2530 3782 2542 3834
rect 2594 3782 2606 3834
rect 2658 3782 19136 3834
rect 1104 3760 19136 3782
rect 2130 3680 2136 3732
rect 2188 3720 2194 3732
rect 2685 3723 2743 3729
rect 2685 3720 2697 3723
rect 2188 3692 2697 3720
rect 2188 3680 2194 3692
rect 2685 3689 2697 3692
rect 2731 3689 2743 3723
rect 2685 3683 2743 3689
rect 6822 3680 6828 3732
rect 6880 3720 6886 3732
rect 7469 3723 7527 3729
rect 7469 3720 7481 3723
rect 6880 3692 7481 3720
rect 6880 3680 6886 3692
rect 7469 3689 7481 3692
rect 7515 3689 7527 3723
rect 7469 3683 7527 3689
rect 10686 3680 10692 3732
rect 10744 3680 10750 3732
rect 11882 3680 11888 3732
rect 11940 3680 11946 3732
rect 12250 3680 12256 3732
rect 12308 3720 12314 3732
rect 12418 3723 12476 3729
rect 12418 3720 12430 3723
rect 12308 3692 12430 3720
rect 12308 3680 12314 3692
rect 12418 3689 12430 3692
rect 12464 3689 12476 3723
rect 12418 3683 12476 3689
rect 12986 3680 12992 3732
rect 13044 3720 13050 3732
rect 13044 3692 15424 3720
rect 13044 3680 13050 3692
rect 6914 3612 6920 3664
rect 6972 3652 6978 3664
rect 15396 3652 15424 3692
rect 15838 3680 15844 3732
rect 15896 3680 15902 3732
rect 15930 3680 15936 3732
rect 15988 3720 15994 3732
rect 16025 3723 16083 3729
rect 16025 3720 16037 3723
rect 15988 3692 16037 3720
rect 15988 3680 15994 3692
rect 16025 3689 16037 3692
rect 16071 3689 16083 3723
rect 16025 3683 16083 3689
rect 17221 3723 17279 3729
rect 17221 3689 17233 3723
rect 17267 3720 17279 3723
rect 17310 3720 17316 3732
rect 17267 3692 17316 3720
rect 17267 3689 17279 3692
rect 17221 3683 17279 3689
rect 17310 3680 17316 3692
rect 17368 3680 17374 3732
rect 18322 3680 18328 3732
rect 18380 3680 18386 3732
rect 18414 3680 18420 3732
rect 18472 3720 18478 3732
rect 18509 3723 18567 3729
rect 18509 3720 18521 3723
rect 18472 3692 18521 3720
rect 18472 3680 18478 3692
rect 18509 3689 18521 3692
rect 18555 3689 18567 3723
rect 18509 3683 18567 3689
rect 17862 3652 17868 3664
rect 6972 3624 8984 3652
rect 15396 3624 17868 3652
rect 6972 3612 6978 3624
rect 2682 3544 2688 3596
rect 2740 3584 2746 3596
rect 5534 3584 5540 3596
rect 2740 3556 5540 3584
rect 2740 3544 2746 3556
rect 5534 3544 5540 3556
rect 5592 3544 5598 3596
rect 5810 3544 5816 3596
rect 5868 3544 5874 3596
rect 7282 3544 7288 3596
rect 7340 3544 7346 3596
rect 8662 3584 8668 3596
rect 7392 3556 8668 3584
rect 842 3476 848 3528
rect 900 3516 906 3528
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 900 3488 1409 3516
rect 900 3476 906 3488
rect 1397 3485 1409 3488
rect 1443 3485 1455 3519
rect 1397 3479 1455 3485
rect 3234 3476 3240 3528
rect 3292 3516 3298 3528
rect 7392 3525 7420 3556
rect 8128 3525 8156 3556
rect 8662 3544 8668 3556
rect 8720 3544 8726 3596
rect 8956 3593 8984 3624
rect 8941 3587 8999 3593
rect 8941 3553 8953 3587
rect 8987 3553 8999 3587
rect 8941 3547 8999 3553
rect 11514 3544 11520 3596
rect 11572 3584 11578 3596
rect 12161 3587 12219 3593
rect 12161 3584 12173 3587
rect 11572 3556 12173 3584
rect 11572 3544 11578 3556
rect 12161 3553 12173 3556
rect 12207 3584 12219 3587
rect 13722 3584 13728 3596
rect 12207 3556 13728 3584
rect 12207 3553 12219 3556
rect 12161 3547 12219 3553
rect 13722 3544 13728 3556
rect 13780 3584 13786 3596
rect 14093 3587 14151 3593
rect 14093 3584 14105 3587
rect 13780 3556 14105 3584
rect 13780 3544 13786 3556
rect 14093 3553 14105 3556
rect 14139 3553 14151 3587
rect 14093 3547 14151 3553
rect 3789 3519 3847 3525
rect 3789 3516 3801 3519
rect 3292 3488 3801 3516
rect 3292 3476 3298 3488
rect 3789 3485 3801 3488
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3485 7435 3519
rect 7377 3479 7435 3485
rect 7561 3519 7619 3525
rect 7561 3485 7573 3519
rect 7607 3485 7619 3519
rect 7561 3479 7619 3485
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3485 8171 3519
rect 8113 3479 8171 3485
rect 7098 3448 7104 3460
rect 7038 3420 7104 3448
rect 7098 3408 7104 3420
rect 7156 3408 7162 3460
rect 7576 3448 7604 3479
rect 8294 3476 8300 3528
rect 8352 3476 8358 3528
rect 8386 3476 8392 3528
rect 8444 3476 8450 3528
rect 8481 3519 8539 3525
rect 8481 3485 8493 3519
rect 8527 3516 8539 3519
rect 8846 3516 8852 3528
rect 8527 3488 8852 3516
rect 8527 3485 8539 3488
rect 8481 3479 8539 3485
rect 8496 3448 8524 3479
rect 8846 3476 8852 3488
rect 8904 3476 8910 3528
rect 11422 3476 11428 3528
rect 11480 3516 11486 3528
rect 11882 3516 11888 3528
rect 11940 3525 11946 3528
rect 11940 3519 11973 3525
rect 11480 3488 11888 3516
rect 11480 3476 11486 3488
rect 11882 3476 11888 3488
rect 11961 3485 11973 3519
rect 11940 3479 11973 3485
rect 12069 3519 12127 3525
rect 12069 3485 12081 3519
rect 12115 3485 12127 3519
rect 12069 3479 12127 3485
rect 11940 3476 11946 3479
rect 7576 3420 8524 3448
rect 8757 3451 8815 3457
rect 3881 3383 3939 3389
rect 3881 3349 3893 3383
rect 3927 3380 3939 3383
rect 3970 3380 3976 3392
rect 3927 3352 3976 3380
rect 3927 3349 3939 3352
rect 3881 3343 3939 3349
rect 3970 3340 3976 3352
rect 4028 3340 4034 3392
rect 6822 3340 6828 3392
rect 6880 3380 6886 3392
rect 7576 3380 7604 3420
rect 8757 3417 8769 3451
rect 8803 3448 8815 3451
rect 9217 3451 9275 3457
rect 9217 3448 9229 3451
rect 8803 3420 9229 3448
rect 8803 3417 8815 3420
rect 8757 3411 8815 3417
rect 9217 3417 9229 3420
rect 9263 3417 9275 3451
rect 9217 3411 9275 3417
rect 9766 3408 9772 3460
rect 9824 3408 9830 3460
rect 6880 3352 7604 3380
rect 12084 3380 12112 3479
rect 13446 3408 13452 3460
rect 13504 3408 13510 3460
rect 13722 3380 13728 3392
rect 12084 3352 13728 3380
rect 6880 3340 6886 3352
rect 13722 3340 13728 3352
rect 13780 3380 13786 3392
rect 13909 3383 13967 3389
rect 13909 3380 13921 3383
rect 13780 3352 13921 3380
rect 13780 3340 13786 3352
rect 13909 3349 13921 3352
rect 13955 3349 13967 3383
rect 14108 3380 14136 3547
rect 15856 3516 15884 3624
rect 17862 3612 17868 3624
rect 17920 3612 17926 3664
rect 17770 3584 17776 3596
rect 17512 3556 17776 3584
rect 15933 3519 15991 3525
rect 15933 3516 15945 3519
rect 15856 3488 15945 3516
rect 15933 3485 15945 3488
rect 15979 3485 15991 3519
rect 15933 3479 15991 3485
rect 16117 3519 16175 3525
rect 16117 3485 16129 3519
rect 16163 3516 16175 3519
rect 16574 3516 16580 3528
rect 16163 3488 16580 3516
rect 16163 3485 16175 3488
rect 16117 3479 16175 3485
rect 16574 3476 16580 3488
rect 16632 3516 16638 3528
rect 17512 3525 17540 3556
rect 17770 3544 17776 3556
rect 17828 3544 17834 3596
rect 18230 3584 18236 3596
rect 18156 3556 18236 3584
rect 17497 3519 17555 3525
rect 17497 3516 17509 3519
rect 16632 3488 17509 3516
rect 16632 3476 16638 3488
rect 17497 3485 17509 3488
rect 17543 3485 17555 3519
rect 17497 3479 17555 3485
rect 17586 3476 17592 3528
rect 17644 3476 17650 3528
rect 17678 3476 17684 3528
rect 17736 3476 17742 3528
rect 17862 3476 17868 3528
rect 17920 3476 17926 3528
rect 18156 3525 18184 3556
rect 18230 3544 18236 3556
rect 18288 3584 18294 3596
rect 18782 3584 18788 3596
rect 18288 3556 18788 3584
rect 18288 3544 18294 3556
rect 18782 3544 18788 3556
rect 18840 3544 18846 3596
rect 18141 3519 18199 3525
rect 18141 3485 18153 3519
rect 18187 3485 18199 3519
rect 18141 3479 18199 3485
rect 18417 3519 18475 3525
rect 18417 3485 18429 3519
rect 18463 3485 18475 3519
rect 18417 3479 18475 3485
rect 14366 3408 14372 3460
rect 14424 3408 14430 3460
rect 15838 3448 15844 3460
rect 15594 3420 15844 3448
rect 15838 3408 15844 3420
rect 15896 3408 15902 3460
rect 16666 3408 16672 3460
rect 16724 3448 16730 3460
rect 17218 3448 17224 3460
rect 16724 3420 17224 3448
rect 16724 3408 16730 3420
rect 17218 3408 17224 3420
rect 17276 3448 17282 3460
rect 18432 3448 18460 3479
rect 17276 3420 18460 3448
rect 17276 3408 17282 3420
rect 17034 3380 17040 3392
rect 14108 3352 17040 3380
rect 13909 3343 13967 3349
rect 17034 3340 17040 3352
rect 17092 3340 17098 3392
rect 1104 3290 19136 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 19136 3290
rect 1104 3216 19136 3238
rect 1581 3179 1639 3185
rect 1581 3145 1593 3179
rect 1627 3176 1639 3179
rect 1670 3176 1676 3188
rect 1627 3148 1676 3176
rect 1627 3145 1639 3148
rect 1581 3139 1639 3145
rect 1670 3136 1676 3148
rect 1728 3136 1734 3188
rect 8754 3176 8760 3188
rect 6472 3148 8760 3176
rect 3970 3068 3976 3120
rect 4028 3068 4034 3120
rect 5629 3111 5687 3117
rect 5629 3108 5641 3111
rect 5198 3080 5641 3108
rect 5629 3077 5641 3080
rect 5675 3077 5687 3111
rect 5629 3071 5687 3077
rect 842 3000 848 3052
rect 900 3040 906 3052
rect 1397 3043 1455 3049
rect 1397 3040 1409 3043
rect 900 3012 1409 3040
rect 900 3000 906 3012
rect 1397 3009 1409 3012
rect 1443 3009 1455 3043
rect 1397 3003 1455 3009
rect 2682 3000 2688 3052
rect 2740 3040 2746 3052
rect 3697 3043 3755 3049
rect 3697 3040 3709 3043
rect 2740 3012 3709 3040
rect 2740 3000 2746 3012
rect 3697 3009 3709 3012
rect 3743 3009 3755 3043
rect 3697 3003 3755 3009
rect 5718 3000 5724 3052
rect 5776 3000 5782 3052
rect 6472 3049 6500 3148
rect 8754 3136 8760 3148
rect 8812 3176 8818 3188
rect 8812 3148 9076 3176
rect 8812 3136 8818 3148
rect 6825 3111 6883 3117
rect 6825 3077 6837 3111
rect 6871 3108 6883 3111
rect 7006 3108 7012 3120
rect 6871 3080 7012 3108
rect 6871 3077 6883 3080
rect 6825 3071 6883 3077
rect 7006 3068 7012 3080
rect 7064 3068 7070 3120
rect 8386 3068 8392 3120
rect 8444 3068 8450 3120
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3009 5871 3043
rect 5813 3003 5871 3009
rect 6457 3043 6515 3049
rect 6457 3009 6469 3043
rect 6503 3009 6515 3043
rect 6457 3003 6515 3009
rect 5445 2975 5503 2981
rect 5445 2941 5457 2975
rect 5491 2972 5503 2975
rect 5828 2972 5856 3003
rect 6914 3000 6920 3052
rect 6972 3040 6978 3052
rect 7101 3043 7159 3049
rect 7101 3040 7113 3043
rect 6972 3012 7113 3040
rect 6972 3000 6978 3012
rect 7101 3009 7113 3012
rect 7147 3009 7159 3043
rect 7101 3003 7159 3009
rect 8941 3043 8999 3049
rect 8941 3009 8953 3043
rect 8987 3009 8999 3043
rect 8941 3003 8999 3009
rect 7377 2975 7435 2981
rect 7377 2972 7389 2975
rect 5491 2944 5856 2972
rect 7024 2944 7389 2972
rect 5491 2941 5503 2944
rect 5445 2935 5503 2941
rect 6638 2864 6644 2916
rect 6696 2904 6702 2916
rect 7024 2913 7052 2944
rect 7377 2941 7389 2944
rect 7423 2941 7435 2975
rect 7377 2935 7435 2941
rect 8849 2975 8907 2981
rect 8849 2941 8861 2975
rect 8895 2972 8907 2975
rect 8956 2972 8984 3003
rect 8895 2944 8984 2972
rect 9048 2972 9076 3148
rect 9766 3136 9772 3188
rect 9824 3136 9830 3188
rect 9858 3136 9864 3188
rect 9916 3176 9922 3188
rect 11698 3176 11704 3188
rect 9916 3148 11704 3176
rect 9916 3136 9922 3148
rect 11698 3136 11704 3148
rect 11756 3136 11762 3188
rect 15194 3136 15200 3188
rect 15252 3176 15258 3188
rect 15657 3179 15715 3185
rect 15657 3176 15669 3179
rect 15252 3148 15669 3176
rect 15252 3136 15258 3148
rect 15657 3145 15669 3148
rect 15703 3145 15715 3179
rect 15657 3139 15715 3145
rect 10873 3111 10931 3117
rect 10873 3077 10885 3111
rect 10919 3108 10931 3111
rect 10962 3108 10968 3120
rect 10919 3080 10968 3108
rect 10919 3077 10931 3080
rect 10873 3071 10931 3077
rect 10962 3068 10968 3080
rect 11020 3068 11026 3120
rect 12066 3108 12072 3120
rect 11072 3080 12072 3108
rect 9677 3043 9735 3049
rect 9677 3009 9689 3043
rect 9723 3040 9735 3043
rect 9858 3040 9864 3052
rect 9723 3012 9864 3040
rect 9723 3009 9735 3012
rect 9677 3003 9735 3009
rect 9858 3000 9864 3012
rect 9916 3000 9922 3052
rect 10045 3043 10103 3049
rect 10045 3009 10057 3043
rect 10091 3040 10103 3043
rect 10686 3040 10692 3052
rect 10091 3012 10692 3040
rect 10091 3009 10103 3012
rect 10045 3003 10103 3009
rect 10686 3000 10692 3012
rect 10744 3000 10750 3052
rect 10505 2975 10563 2981
rect 10505 2972 10517 2975
rect 9048 2944 10517 2972
rect 8895 2941 8907 2944
rect 8849 2935 8907 2941
rect 10505 2941 10517 2944
rect 10551 2972 10563 2975
rect 11072 2972 11100 3080
rect 12066 3068 12072 3080
rect 12124 3068 12130 3120
rect 12526 3068 12532 3120
rect 12584 3068 12590 3120
rect 15470 3068 15476 3120
rect 15528 3068 15534 3120
rect 15672 3108 15700 3139
rect 15838 3136 15844 3188
rect 15896 3136 15902 3188
rect 16942 3176 16948 3188
rect 16546 3148 16948 3176
rect 16546 3108 16574 3148
rect 16942 3136 16948 3148
rect 17000 3136 17006 3188
rect 17034 3108 17040 3120
rect 15672 3080 16574 3108
rect 16684 3080 17040 3108
rect 11141 3043 11199 3049
rect 11141 3009 11153 3043
rect 11187 3040 11199 3043
rect 11238 3040 11244 3052
rect 11187 3012 11244 3040
rect 11187 3009 11199 3012
rect 11141 3003 11199 3009
rect 11238 3000 11244 3012
rect 11296 3000 11302 3052
rect 11514 3000 11520 3052
rect 11572 3000 11578 3052
rect 13357 3043 13415 3049
rect 13357 3040 13369 3043
rect 13280 3012 13369 3040
rect 11793 2975 11851 2981
rect 11793 2972 11805 2975
rect 10551 2944 11100 2972
rect 11164 2944 11805 2972
rect 10551 2941 10563 2944
rect 10505 2935 10563 2941
rect 11164 2916 11192 2944
rect 11793 2941 11805 2944
rect 11839 2941 11851 2975
rect 11793 2935 11851 2941
rect 11882 2932 11888 2984
rect 11940 2972 11946 2984
rect 12434 2972 12440 2984
rect 11940 2944 12440 2972
rect 11940 2932 11946 2944
rect 12434 2932 12440 2944
rect 12492 2932 12498 2984
rect 13280 2981 13308 3012
rect 13357 3009 13369 3012
rect 13403 3009 13415 3043
rect 13357 3003 13415 3009
rect 13722 3000 13728 3052
rect 13780 3000 13786 3052
rect 16684 3049 16712 3080
rect 17034 3068 17040 3080
rect 17092 3068 17098 3120
rect 17218 3068 17224 3120
rect 17276 3108 17282 3120
rect 17276 3080 17434 3108
rect 17276 3068 17282 3080
rect 15933 3043 15991 3049
rect 15933 3009 15945 3043
rect 15979 3040 15991 3043
rect 16658 3043 16716 3049
rect 15979 3012 16574 3040
rect 15979 3009 15991 3012
rect 15933 3003 15991 3009
rect 13265 2975 13323 2981
rect 13265 2941 13277 2975
rect 13311 2941 13323 2975
rect 13265 2935 13323 2941
rect 15105 2975 15163 2981
rect 15105 2941 15117 2975
rect 15151 2972 15163 2975
rect 16022 2972 16028 2984
rect 15151 2944 16028 2972
rect 15151 2941 15163 2944
rect 15105 2935 15163 2941
rect 7009 2907 7067 2913
rect 7009 2904 7021 2907
rect 6696 2876 7021 2904
rect 6696 2864 6702 2876
rect 7009 2873 7021 2876
rect 7055 2873 7067 2907
rect 7009 2867 7067 2873
rect 11057 2907 11115 2913
rect 11057 2873 11069 2907
rect 11103 2904 11115 2907
rect 11146 2904 11152 2916
rect 11103 2876 11152 2904
rect 11103 2873 11115 2876
rect 11057 2867 11115 2873
rect 11146 2864 11152 2876
rect 11204 2864 11210 2916
rect 11422 2904 11428 2916
rect 11256 2876 11428 2904
rect 5997 2839 6055 2845
rect 5997 2805 6009 2839
rect 6043 2836 6055 2839
rect 6730 2836 6736 2848
rect 6043 2808 6736 2836
rect 6043 2805 6055 2808
rect 5997 2799 6055 2805
rect 6730 2796 6736 2808
rect 6788 2796 6794 2848
rect 6822 2796 6828 2848
rect 6880 2796 6886 2848
rect 9125 2839 9183 2845
rect 9125 2805 9137 2839
rect 9171 2836 9183 2839
rect 9306 2836 9312 2848
rect 9171 2808 9312 2836
rect 9171 2805 9183 2808
rect 9125 2799 9183 2805
rect 9306 2796 9312 2808
rect 9364 2796 9370 2848
rect 10229 2839 10287 2845
rect 10229 2805 10241 2839
rect 10275 2836 10287 2839
rect 10594 2836 10600 2848
rect 10275 2808 10600 2836
rect 10275 2805 10287 2808
rect 10229 2799 10287 2805
rect 10594 2796 10600 2808
rect 10652 2796 10658 2848
rect 10873 2839 10931 2845
rect 10873 2805 10885 2839
rect 10919 2836 10931 2839
rect 11256 2836 11284 2876
rect 11422 2864 11428 2876
rect 11480 2864 11486 2916
rect 15120 2904 15148 2935
rect 16022 2932 16028 2944
rect 16080 2932 16086 2984
rect 16546 2904 16574 3012
rect 16658 3009 16670 3043
rect 16704 3009 16716 3043
rect 16658 3003 16716 3009
rect 18509 3043 18567 3049
rect 18509 3009 18521 3043
rect 18555 3009 18567 3043
rect 18509 3003 18567 3009
rect 16942 2932 16948 2984
rect 17000 2932 17006 2984
rect 18417 2975 18475 2981
rect 18417 2941 18429 2975
rect 18463 2972 18475 2975
rect 18524 2972 18552 3003
rect 18463 2944 18552 2972
rect 18463 2941 18475 2944
rect 18417 2935 18475 2941
rect 16666 2904 16672 2916
rect 12820 2876 15148 2904
rect 15488 2876 16068 2904
rect 16546 2876 16672 2904
rect 10919 2808 11284 2836
rect 11333 2839 11391 2845
rect 10919 2805 10931 2808
rect 10873 2799 10931 2805
rect 11333 2805 11345 2839
rect 11379 2836 11391 2839
rect 12158 2836 12164 2848
rect 11379 2808 12164 2836
rect 11379 2805 11391 2808
rect 11333 2799 11391 2805
rect 12158 2796 12164 2808
rect 12216 2796 12222 2848
rect 12250 2796 12256 2848
rect 12308 2836 12314 2848
rect 12820 2836 12848 2876
rect 12308 2808 12848 2836
rect 13541 2839 13599 2845
rect 12308 2796 12314 2808
rect 13541 2805 13553 2839
rect 13587 2836 13599 2839
rect 13814 2836 13820 2848
rect 13587 2808 13820 2836
rect 13587 2805 13599 2808
rect 13541 2799 13599 2805
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 13909 2839 13967 2845
rect 13909 2805 13921 2839
rect 13955 2836 13967 2839
rect 14458 2836 14464 2848
rect 13955 2808 14464 2836
rect 13955 2805 13967 2808
rect 13909 2799 13967 2805
rect 14458 2796 14464 2808
rect 14516 2796 14522 2848
rect 15488 2845 15516 2876
rect 15473 2839 15531 2845
rect 15473 2805 15485 2839
rect 15519 2805 15531 2839
rect 16040 2836 16068 2876
rect 16666 2864 16672 2876
rect 16724 2864 16730 2916
rect 16574 2836 16580 2848
rect 16040 2808 16580 2836
rect 15473 2799 15531 2805
rect 16574 2796 16580 2808
rect 16632 2796 16638 2848
rect 18598 2796 18604 2848
rect 18656 2836 18662 2848
rect 18693 2839 18751 2845
rect 18693 2836 18705 2839
rect 18656 2808 18705 2836
rect 18656 2796 18662 2808
rect 18693 2805 18705 2808
rect 18739 2805 18751 2839
rect 18693 2799 18751 2805
rect 1104 2746 19136 2768
rect 1104 2694 2350 2746
rect 2402 2694 2414 2746
rect 2466 2694 2478 2746
rect 2530 2694 2542 2746
rect 2594 2694 2606 2746
rect 2658 2694 19136 2746
rect 1104 2672 19136 2694
rect 6089 2635 6147 2641
rect 6089 2601 6101 2635
rect 6135 2632 6147 2635
rect 6822 2632 6828 2644
rect 6135 2604 6828 2632
rect 6135 2601 6147 2604
rect 6089 2595 6147 2601
rect 6822 2592 6828 2604
rect 6880 2592 6886 2644
rect 7006 2592 7012 2644
rect 7064 2632 7070 2644
rect 7193 2635 7251 2641
rect 7193 2632 7205 2635
rect 7064 2604 7205 2632
rect 7064 2592 7070 2604
rect 7193 2601 7205 2604
rect 7239 2601 7251 2635
rect 7193 2595 7251 2601
rect 8205 2635 8263 2641
rect 8205 2601 8217 2635
rect 8251 2632 8263 2635
rect 8386 2632 8392 2644
rect 8251 2604 8392 2632
rect 8251 2601 8263 2604
rect 8205 2595 8263 2601
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 11054 2592 11060 2644
rect 11112 2592 11118 2644
rect 11793 2635 11851 2641
rect 11793 2601 11805 2635
rect 11839 2632 11851 2635
rect 12526 2632 12532 2644
rect 11839 2604 12532 2632
rect 11839 2601 11851 2604
rect 11793 2595 11851 2601
rect 12526 2592 12532 2604
rect 12584 2592 12590 2644
rect 15470 2592 15476 2644
rect 15528 2632 15534 2644
rect 15565 2635 15623 2641
rect 15565 2632 15577 2635
rect 15528 2604 15577 2632
rect 15528 2592 15534 2604
rect 15565 2601 15577 2604
rect 15611 2601 15623 2635
rect 15565 2595 15623 2601
rect 17218 2592 17224 2644
rect 17276 2632 17282 2644
rect 17313 2635 17371 2641
rect 17313 2632 17325 2635
rect 17276 2604 17325 2632
rect 17276 2592 17282 2604
rect 17313 2601 17325 2604
rect 17359 2601 17371 2635
rect 17313 2595 17371 2601
rect 17402 2592 17408 2644
rect 17460 2632 17466 2644
rect 17497 2635 17555 2641
rect 17497 2632 17509 2635
rect 17460 2604 17509 2632
rect 17460 2592 17466 2604
rect 17497 2601 17509 2604
rect 17543 2601 17555 2635
rect 17497 2595 17555 2601
rect 17770 2592 17776 2644
rect 17828 2592 17834 2644
rect 18046 2592 18052 2644
rect 18104 2592 18110 2644
rect 18782 2592 18788 2644
rect 18840 2592 18846 2644
rect 8021 2567 8079 2573
rect 8021 2533 8033 2567
rect 8067 2564 8079 2567
rect 8570 2564 8576 2576
rect 8067 2536 8576 2564
rect 8067 2533 8079 2536
rect 8021 2527 8079 2533
rect 8570 2524 8576 2536
rect 8628 2524 8634 2576
rect 11606 2524 11612 2576
rect 11664 2564 11670 2576
rect 11977 2567 12035 2573
rect 11977 2564 11989 2567
rect 11664 2536 11989 2564
rect 11664 2524 11670 2536
rect 11977 2533 11989 2536
rect 12023 2533 12035 2567
rect 11977 2527 12035 2533
rect 16482 2524 16488 2576
rect 16540 2564 16546 2576
rect 18325 2567 18383 2573
rect 18325 2564 18337 2567
rect 16540 2536 18337 2564
rect 16540 2524 16546 2536
rect 18325 2533 18337 2536
rect 18371 2533 18383 2567
rect 18325 2527 18383 2533
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 5868 2400 5917 2428
rect 5868 2388 5874 2400
rect 5905 2397 5917 2400
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 6730 2388 6736 2440
rect 6788 2388 6794 2440
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7377 2431 7435 2437
rect 7377 2428 7389 2431
rect 7156 2400 7389 2428
rect 7156 2388 7162 2400
rect 7377 2397 7389 2400
rect 7423 2397 7435 2431
rect 7377 2391 7435 2397
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 7837 2431 7895 2437
rect 7837 2428 7849 2431
rect 7800 2400 7849 2428
rect 7800 2388 7806 2400
rect 7837 2397 7849 2400
rect 7883 2397 7895 2431
rect 7837 2391 7895 2397
rect 8110 2388 8116 2440
rect 8168 2388 8174 2440
rect 9306 2388 9312 2440
rect 9364 2388 9370 2440
rect 10594 2388 10600 2440
rect 10652 2388 10658 2440
rect 10962 2388 10968 2440
rect 11020 2428 11026 2440
rect 11241 2431 11299 2437
rect 11241 2428 11253 2431
rect 11020 2400 11253 2428
rect 11020 2388 11026 2400
rect 11241 2397 11253 2400
rect 11287 2397 11299 2431
rect 11241 2391 11299 2397
rect 11698 2388 11704 2440
rect 11756 2388 11762 2440
rect 12158 2388 12164 2440
rect 12216 2388 12222 2440
rect 12250 2388 12256 2440
rect 12308 2428 12314 2440
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 12308 2400 12357 2428
rect 12308 2388 12314 2400
rect 12345 2397 12357 2400
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 13814 2388 13820 2440
rect 13872 2388 13878 2440
rect 14458 2388 14464 2440
rect 14516 2388 14522 2440
rect 15470 2388 15476 2440
rect 15528 2428 15534 2440
rect 15749 2431 15807 2437
rect 15749 2428 15761 2431
rect 15528 2400 15761 2428
rect 15528 2388 15534 2400
rect 15749 2397 15761 2400
rect 15795 2397 15807 2431
rect 15749 2391 15807 2397
rect 16666 2388 16672 2440
rect 16724 2428 16730 2440
rect 17221 2431 17279 2437
rect 17221 2428 17233 2431
rect 16724 2400 17233 2428
rect 16724 2388 16730 2400
rect 17221 2397 17233 2400
rect 17267 2397 17279 2431
rect 17221 2391 17279 2397
rect 17678 2388 17684 2440
rect 17736 2388 17742 2440
rect 17954 2388 17960 2440
rect 18012 2388 18018 2440
rect 18230 2388 18236 2440
rect 18288 2388 18294 2440
rect 18506 2388 18512 2440
rect 18564 2388 18570 2440
rect 18598 2388 18604 2440
rect 18656 2388 18662 2440
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6549 2295 6607 2301
rect 6549 2292 6561 2295
rect 6512 2264 6561 2292
rect 6512 2252 6518 2264
rect 6549 2261 6561 2264
rect 6595 2261 6607 2295
rect 6549 2255 6607 2261
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 9125 2295 9183 2301
rect 9125 2292 9137 2295
rect 9088 2264 9137 2292
rect 9088 2252 9094 2264
rect 9125 2261 9137 2264
rect 9171 2261 9183 2295
rect 9125 2255 9183 2261
rect 10318 2252 10324 2304
rect 10376 2292 10382 2304
rect 10413 2295 10471 2301
rect 10413 2292 10425 2295
rect 10376 2264 10425 2292
rect 10376 2252 10382 2264
rect 10413 2261 10425 2264
rect 10459 2261 10471 2295
rect 10413 2255 10471 2261
rect 12434 2252 12440 2304
rect 12492 2292 12498 2304
rect 12529 2295 12587 2301
rect 12529 2292 12541 2295
rect 12492 2264 12541 2292
rect 12492 2252 12498 2264
rect 12529 2261 12541 2264
rect 12575 2261 12587 2295
rect 12529 2255 12587 2261
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 13633 2295 13691 2301
rect 13633 2292 13645 2295
rect 13596 2264 13645 2292
rect 13596 2252 13602 2264
rect 13633 2261 13645 2264
rect 13679 2261 13691 2295
rect 13633 2255 13691 2261
rect 14182 2252 14188 2304
rect 14240 2292 14246 2304
rect 14277 2295 14335 2301
rect 14277 2292 14289 2295
rect 14240 2264 14289 2292
rect 14240 2252 14246 2264
rect 14277 2261 14289 2264
rect 14323 2261 14335 2295
rect 14277 2255 14335 2261
rect 1104 2202 19136 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 19136 2202
rect 1104 2128 19136 2150
<< via1 >>
rect 2350 20102 2402 20154
rect 2414 20102 2466 20154
rect 2478 20102 2530 20154
rect 2542 20102 2594 20154
rect 2606 20102 2658 20154
rect 5264 20043 5316 20052
rect 5264 20009 5273 20043
rect 5273 20009 5307 20043
rect 5307 20009 5316 20043
rect 5264 20000 5316 20009
rect 8484 20043 8536 20052
rect 8484 20009 8493 20043
rect 8493 20009 8527 20043
rect 8527 20009 8536 20043
rect 8484 20000 8536 20009
rect 9772 20043 9824 20052
rect 9772 20009 9781 20043
rect 9781 20009 9815 20043
rect 9815 20009 9824 20043
rect 9772 20000 9824 20009
rect 10876 20000 10928 20052
rect 11704 20043 11756 20052
rect 11704 20009 11713 20043
rect 11713 20009 11747 20043
rect 11747 20009 11756 20043
rect 11704 20000 11756 20009
rect 12992 20043 13044 20052
rect 12992 20009 13001 20043
rect 13001 20009 13035 20043
rect 13035 20009 13044 20043
rect 12992 20000 13044 20009
rect 14280 20043 14332 20052
rect 14280 20009 14289 20043
rect 14289 20009 14323 20043
rect 14323 20009 14332 20043
rect 14280 20000 14332 20009
rect 17500 20043 17552 20052
rect 17500 20009 17509 20043
rect 17509 20009 17543 20043
rect 17543 20009 17552 20043
rect 17500 20000 17552 20009
rect 17776 20043 17828 20052
rect 17776 20009 17785 20043
rect 17785 20009 17819 20043
rect 17819 20009 17828 20043
rect 17776 20000 17828 20009
rect 4896 19796 4948 19848
rect 5908 19839 5960 19848
rect 5908 19805 5917 19839
rect 5917 19805 5951 19839
rect 5951 19805 5960 19839
rect 5908 19796 5960 19805
rect 6736 19839 6788 19848
rect 6736 19805 6745 19839
rect 6745 19805 6779 19839
rect 6779 19805 6788 19839
rect 6736 19796 6788 19805
rect 7196 19839 7248 19848
rect 7196 19805 7205 19839
rect 7205 19805 7239 19839
rect 7239 19805 7248 19839
rect 7196 19796 7248 19805
rect 8668 19839 8720 19848
rect 8668 19805 8677 19839
rect 8677 19805 8711 19839
rect 8711 19805 8720 19839
rect 8668 19796 8720 19805
rect 9956 19839 10008 19848
rect 9956 19805 9965 19839
rect 9965 19805 9999 19839
rect 9999 19805 10008 19839
rect 9956 19796 10008 19805
rect 9496 19728 9548 19780
rect 10600 19796 10652 19848
rect 11704 19796 11756 19848
rect 13268 19796 13320 19848
rect 13728 19796 13780 19848
rect 14464 19839 14516 19848
rect 14464 19805 14473 19839
rect 14473 19805 14507 19839
rect 14507 19805 14516 19839
rect 14464 19796 14516 19805
rect 14924 19839 14976 19848
rect 14924 19805 14933 19839
rect 14933 19805 14967 19839
rect 14967 19805 14976 19839
rect 14924 19796 14976 19805
rect 16212 19839 16264 19848
rect 16212 19805 16221 19839
rect 16221 19805 16255 19839
rect 16255 19805 16264 19839
rect 16212 19796 16264 19805
rect 17868 19839 17920 19848
rect 17868 19805 17877 19839
rect 17877 19805 17911 19839
rect 17911 19805 17920 19839
rect 17868 19796 17920 19805
rect 18236 19796 18288 19848
rect 18512 19796 18564 19848
rect 5724 19660 5776 19712
rect 6552 19703 6604 19712
rect 6552 19669 6561 19703
rect 6561 19669 6595 19703
rect 6595 19669 6604 19703
rect 6552 19660 6604 19669
rect 8392 19660 8444 19712
rect 9404 19660 9456 19712
rect 10508 19660 10560 19712
rect 12900 19660 12952 19712
rect 14924 19660 14976 19712
rect 16396 19703 16448 19712
rect 16396 19669 16405 19703
rect 16405 19669 16439 19703
rect 16439 19669 16448 19703
rect 16396 19660 16448 19669
rect 18052 19703 18104 19712
rect 18052 19669 18061 19703
rect 18061 19669 18095 19703
rect 18095 19669 18104 19703
rect 18052 19660 18104 19669
rect 3010 19558 3062 19610
rect 3074 19558 3126 19610
rect 3138 19558 3190 19610
rect 3202 19558 3254 19610
rect 3266 19558 3318 19610
rect 2872 19388 2924 19440
rect 3976 19388 4028 19440
rect 4896 19499 4948 19508
rect 4896 19465 4905 19499
rect 4905 19465 4939 19499
rect 4939 19465 4948 19499
rect 4896 19456 4948 19465
rect 6552 19499 6604 19508
rect 6552 19465 6561 19499
rect 6561 19465 6595 19499
rect 6595 19465 6604 19499
rect 6552 19456 6604 19465
rect 9496 19499 9548 19508
rect 9496 19465 9505 19499
rect 9505 19465 9539 19499
rect 9539 19465 9548 19499
rect 9496 19456 9548 19465
rect 5724 19363 5776 19372
rect 5724 19329 5733 19363
rect 5733 19329 5767 19363
rect 5767 19329 5776 19363
rect 5724 19320 5776 19329
rect 5908 19363 5960 19372
rect 5908 19329 5917 19363
rect 5917 19329 5951 19363
rect 5951 19329 5960 19363
rect 5908 19320 5960 19329
rect 6644 19388 6696 19440
rect 6736 19320 6788 19372
rect 9312 19388 9364 19440
rect 11704 19499 11756 19508
rect 11704 19465 11713 19499
rect 11713 19465 11747 19499
rect 11747 19465 11756 19499
rect 11704 19456 11756 19465
rect 13268 19499 13320 19508
rect 13268 19465 13277 19499
rect 13277 19465 13311 19499
rect 13311 19465 13320 19499
rect 13268 19456 13320 19465
rect 14464 19456 14516 19508
rect 14924 19499 14976 19508
rect 14924 19465 14933 19499
rect 14933 19465 14967 19499
rect 14967 19465 14976 19499
rect 14924 19456 14976 19465
rect 17868 19456 17920 19508
rect 9588 19363 9640 19372
rect 9588 19329 9597 19363
rect 9597 19329 9631 19363
rect 9631 19329 9640 19363
rect 9588 19320 9640 19329
rect 10968 19320 11020 19372
rect 11520 19363 11572 19372
rect 11520 19329 11529 19363
rect 11529 19329 11563 19363
rect 11563 19329 11572 19363
rect 11520 19320 11572 19329
rect 12900 19363 12952 19372
rect 12900 19329 12908 19363
rect 12908 19329 12942 19363
rect 12942 19329 12952 19363
rect 12900 19320 12952 19329
rect 16948 19388 17000 19440
rect 8760 19252 8812 19304
rect 10600 19252 10652 19304
rect 13636 19363 13688 19372
rect 13636 19329 13645 19363
rect 13645 19329 13679 19363
rect 13679 19329 13688 19363
rect 13636 19320 13688 19329
rect 15200 19363 15252 19372
rect 15200 19329 15209 19363
rect 15209 19329 15243 19363
rect 15243 19329 15252 19363
rect 15200 19320 15252 19329
rect 16396 19320 16448 19372
rect 18696 19363 18748 19372
rect 18696 19329 18705 19363
rect 18705 19329 18739 19363
rect 18739 19329 18748 19363
rect 18696 19320 18748 19329
rect 2688 19184 2740 19236
rect 5724 19184 5776 19236
rect 5632 19116 5684 19168
rect 5816 19159 5868 19168
rect 5816 19125 5825 19159
rect 5825 19125 5859 19159
rect 5859 19125 5868 19159
rect 5816 19116 5868 19125
rect 6460 19116 6512 19168
rect 6828 19116 6880 19168
rect 7196 19116 7248 19168
rect 10232 19116 10284 19168
rect 11796 19116 11848 19168
rect 12716 19116 12768 19168
rect 16672 19295 16724 19304
rect 16672 19261 16681 19295
rect 16681 19261 16715 19295
rect 16715 19261 16724 19295
rect 16672 19252 16724 19261
rect 14832 19184 14884 19236
rect 15292 19159 15344 19168
rect 15292 19125 15301 19159
rect 15301 19125 15335 19159
rect 15335 19125 15344 19159
rect 15292 19116 15344 19125
rect 18420 19159 18472 19168
rect 18420 19125 18429 19159
rect 18429 19125 18463 19159
rect 18463 19125 18472 19159
rect 18420 19116 18472 19125
rect 2350 19014 2402 19066
rect 2414 19014 2466 19066
rect 2478 19014 2530 19066
rect 2542 19014 2594 19066
rect 2606 19014 2658 19066
rect 3976 18912 4028 18964
rect 8668 18912 8720 18964
rect 8760 18912 8812 18964
rect 9312 18912 9364 18964
rect 10232 18844 10284 18896
rect 10600 18912 10652 18964
rect 10968 18912 11020 18964
rect 13636 18912 13688 18964
rect 16948 18955 17000 18964
rect 16948 18921 16957 18955
rect 16957 18921 16991 18955
rect 16991 18921 17000 18955
rect 16948 18912 17000 18921
rect 18052 18955 18104 18964
rect 18052 18921 18061 18955
rect 18061 18921 18095 18955
rect 18095 18921 18104 18955
rect 18052 18912 18104 18921
rect 11704 18844 11756 18896
rect 848 18708 900 18760
rect 1676 18708 1728 18760
rect 6552 18776 6604 18828
rect 3976 18751 4028 18760
rect 3976 18717 3985 18751
rect 3985 18717 4019 18751
rect 4019 18717 4028 18751
rect 3976 18708 4028 18717
rect 9128 18776 9180 18828
rect 8392 18708 8444 18760
rect 9680 18776 9732 18828
rect 9404 18751 9456 18760
rect 9404 18717 9413 18751
rect 9413 18717 9447 18751
rect 9447 18717 9456 18751
rect 9404 18708 9456 18717
rect 11152 18776 11204 18828
rect 12624 18776 12676 18828
rect 2320 18640 2372 18692
rect 3424 18640 3476 18692
rect 4620 18683 4672 18692
rect 4620 18649 4629 18683
rect 4629 18649 4663 18683
rect 4663 18649 4672 18683
rect 4620 18640 4672 18649
rect 5632 18640 5684 18692
rect 6460 18683 6512 18692
rect 6460 18649 6469 18683
rect 6469 18649 6503 18683
rect 6503 18649 6512 18683
rect 6460 18640 6512 18649
rect 7196 18640 7248 18692
rect 1768 18572 1820 18624
rect 3516 18615 3568 18624
rect 3516 18581 3525 18615
rect 3525 18581 3559 18615
rect 3559 18581 3568 18615
rect 3516 18572 3568 18581
rect 6000 18572 6052 18624
rect 7380 18572 7432 18624
rect 16396 18708 16448 18760
rect 10508 18683 10560 18692
rect 10508 18649 10517 18683
rect 10517 18649 10551 18683
rect 10551 18649 10560 18683
rect 10508 18640 10560 18649
rect 12164 18640 12216 18692
rect 12992 18640 13044 18692
rect 14648 18640 14700 18692
rect 15384 18640 15436 18692
rect 16856 18751 16908 18760
rect 16856 18717 16865 18751
rect 16865 18717 16899 18751
rect 16899 18717 16908 18751
rect 16856 18708 16908 18717
rect 18328 18751 18380 18760
rect 18328 18717 18337 18751
rect 18337 18717 18371 18751
rect 18371 18717 18380 18751
rect 18328 18708 18380 18717
rect 18420 18751 18472 18760
rect 18420 18717 18429 18751
rect 18429 18717 18463 18751
rect 18463 18717 18472 18751
rect 18420 18708 18472 18717
rect 11428 18572 11480 18624
rect 15660 18572 15712 18624
rect 16488 18572 16540 18624
rect 18604 18615 18656 18624
rect 18604 18581 18613 18615
rect 18613 18581 18647 18615
rect 18647 18581 18656 18615
rect 18604 18572 18656 18581
rect 3010 18470 3062 18522
rect 3074 18470 3126 18522
rect 3138 18470 3190 18522
rect 3202 18470 3254 18522
rect 3266 18470 3318 18522
rect 1768 18411 1820 18420
rect 1768 18377 1777 18411
rect 1777 18377 1811 18411
rect 1811 18377 1820 18411
rect 1768 18368 1820 18377
rect 2320 18411 2372 18420
rect 2320 18377 2329 18411
rect 2329 18377 2363 18411
rect 2363 18377 2372 18411
rect 2320 18368 2372 18377
rect 3424 18368 3476 18420
rect 4620 18368 4672 18420
rect 5816 18368 5868 18420
rect 6828 18368 6880 18420
rect 2596 18300 2648 18352
rect 2688 18232 2740 18284
rect 2964 18232 3016 18284
rect 3332 18275 3384 18284
rect 3332 18241 3341 18275
rect 3341 18241 3375 18275
rect 3375 18241 3384 18275
rect 3332 18232 3384 18241
rect 3976 18232 4028 18284
rect 6460 18300 6512 18352
rect 6000 18275 6052 18284
rect 6000 18241 6009 18275
rect 6009 18241 6043 18275
rect 6043 18241 6052 18275
rect 6000 18232 6052 18241
rect 3516 18164 3568 18216
rect 5908 18164 5960 18216
rect 7380 18232 7432 18284
rect 6736 18207 6788 18216
rect 6736 18173 6745 18207
rect 6745 18173 6779 18207
rect 6779 18173 6788 18207
rect 6736 18164 6788 18173
rect 7564 18275 7616 18284
rect 7564 18241 7573 18275
rect 7573 18241 7607 18275
rect 7607 18241 7616 18275
rect 7564 18232 7616 18241
rect 9956 18368 10008 18420
rect 12164 18411 12216 18420
rect 12164 18377 12173 18411
rect 12173 18377 12207 18411
rect 12207 18377 12216 18411
rect 12164 18368 12216 18377
rect 11428 18300 11480 18352
rect 9220 18275 9272 18284
rect 9220 18241 9229 18275
rect 9229 18241 9263 18275
rect 9263 18241 9272 18275
rect 9220 18232 9272 18241
rect 12532 18281 12584 18308
rect 12532 18256 12538 18281
rect 12538 18256 12572 18281
rect 12572 18256 12584 18281
rect 11704 18164 11756 18216
rect 12716 18232 12768 18284
rect 12992 18368 13044 18420
rect 14648 18411 14700 18420
rect 14648 18377 14657 18411
rect 14657 18377 14691 18411
rect 14691 18377 14700 18411
rect 14648 18368 14700 18377
rect 15292 18368 15344 18420
rect 18328 18368 18380 18420
rect 18788 18411 18840 18420
rect 18788 18377 18797 18411
rect 18797 18377 18831 18411
rect 18831 18377 18840 18411
rect 18788 18368 18840 18377
rect 12900 18164 12952 18216
rect 1952 18096 2004 18148
rect 2780 18096 2832 18148
rect 3332 18096 3384 18148
rect 11152 18096 11204 18148
rect 12716 18096 12768 18148
rect 14832 18275 14884 18284
rect 14832 18241 14841 18275
rect 14841 18241 14875 18275
rect 14875 18241 14884 18275
rect 14832 18232 14884 18241
rect 17684 18300 17736 18352
rect 15660 18232 15712 18284
rect 18604 18275 18656 18284
rect 18604 18241 18613 18275
rect 18613 18241 18647 18275
rect 18647 18241 18656 18275
rect 18604 18232 18656 18241
rect 15752 18207 15804 18216
rect 15752 18173 15761 18207
rect 15761 18173 15795 18207
rect 15795 18173 15804 18207
rect 15752 18164 15804 18173
rect 15844 18164 15896 18216
rect 16672 18207 16724 18216
rect 16672 18173 16681 18207
rect 16681 18173 16715 18207
rect 16715 18173 16724 18207
rect 16672 18164 16724 18173
rect 16948 18207 17000 18216
rect 16948 18173 16957 18207
rect 16957 18173 16991 18207
rect 16991 18173 17000 18207
rect 16948 18164 17000 18173
rect 15384 18096 15436 18148
rect 1584 18028 1636 18080
rect 2228 18028 2280 18080
rect 2596 18028 2648 18080
rect 2964 18028 3016 18080
rect 3424 18028 3476 18080
rect 5908 18028 5960 18080
rect 7932 18071 7984 18080
rect 7932 18037 7941 18071
rect 7941 18037 7975 18071
rect 7975 18037 7984 18071
rect 7932 18028 7984 18037
rect 16580 18028 16632 18080
rect 2350 17926 2402 17978
rect 2414 17926 2466 17978
rect 2478 17926 2530 17978
rect 2542 17926 2594 17978
rect 2606 17926 2658 17978
rect 1584 17867 1636 17876
rect 1584 17833 1593 17867
rect 1593 17833 1627 17867
rect 1627 17833 1636 17867
rect 1584 17824 1636 17833
rect 12348 17867 12400 17876
rect 12348 17833 12357 17867
rect 12357 17833 12391 17867
rect 12391 17833 12400 17867
rect 12348 17824 12400 17833
rect 16948 17867 17000 17876
rect 16948 17833 16957 17867
rect 16957 17833 16991 17867
rect 16991 17833 17000 17867
rect 16948 17824 17000 17833
rect 17684 17867 17736 17876
rect 17684 17833 17693 17867
rect 17693 17833 17727 17867
rect 17727 17833 17736 17867
rect 17684 17824 17736 17833
rect 6736 17799 6788 17808
rect 6736 17765 6745 17799
rect 6745 17765 6779 17799
rect 6779 17765 6788 17799
rect 6736 17756 6788 17765
rect 848 17620 900 17672
rect 6368 17663 6420 17672
rect 6368 17629 6377 17663
rect 6377 17629 6411 17663
rect 6411 17629 6420 17663
rect 6368 17620 6420 17629
rect 6460 17663 6512 17672
rect 6460 17629 6470 17663
rect 6470 17629 6504 17663
rect 6504 17629 6512 17663
rect 6460 17620 6512 17629
rect 8668 17620 8720 17672
rect 10600 17663 10652 17672
rect 10600 17629 10609 17663
rect 10609 17629 10643 17663
rect 10643 17629 10652 17663
rect 10600 17620 10652 17629
rect 11336 17688 11388 17740
rect 16396 17688 16448 17740
rect 11152 17663 11204 17672
rect 11152 17629 11161 17663
rect 11161 17629 11195 17663
rect 11195 17629 11204 17663
rect 11152 17620 11204 17629
rect 11888 17620 11940 17672
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 14832 17552 14884 17604
rect 15292 17552 15344 17604
rect 16488 17663 16540 17672
rect 16488 17629 16497 17663
rect 16497 17629 16531 17663
rect 16531 17629 16540 17663
rect 16488 17620 16540 17629
rect 16580 17663 16632 17672
rect 16580 17629 16589 17663
rect 16589 17629 16623 17663
rect 16623 17629 16632 17663
rect 16580 17620 16632 17629
rect 16856 17620 16908 17672
rect 17868 17620 17920 17672
rect 18788 17663 18840 17672
rect 18788 17629 18797 17663
rect 18797 17629 18831 17663
rect 18831 17629 18840 17663
rect 18788 17620 18840 17629
rect 17776 17552 17828 17604
rect 8576 17484 8628 17536
rect 9864 17484 9916 17536
rect 10784 17527 10836 17536
rect 10784 17493 10793 17527
rect 10793 17493 10827 17527
rect 10827 17493 10836 17527
rect 10784 17484 10836 17493
rect 10876 17484 10928 17536
rect 15200 17484 15252 17536
rect 18144 17484 18196 17536
rect 3010 17382 3062 17434
rect 3074 17382 3126 17434
rect 3138 17382 3190 17434
rect 3202 17382 3254 17434
rect 3266 17382 3318 17434
rect 9220 17280 9272 17332
rect 10784 17280 10836 17332
rect 11888 17323 11940 17332
rect 11888 17289 11897 17323
rect 11897 17289 11931 17323
rect 11931 17289 11940 17323
rect 11888 17280 11940 17289
rect 14832 17280 14884 17332
rect 15752 17280 15804 17332
rect 1216 17212 1268 17264
rect 1584 17187 1636 17196
rect 1584 17153 1593 17187
rect 1593 17153 1627 17187
rect 1627 17153 1636 17187
rect 1584 17144 1636 17153
rect 2136 17144 2188 17196
rect 2320 17187 2372 17196
rect 2320 17153 2329 17187
rect 2329 17153 2363 17187
rect 2363 17153 2372 17187
rect 2320 17144 2372 17153
rect 6552 17255 6604 17264
rect 6552 17221 6561 17255
rect 6561 17221 6595 17255
rect 6595 17221 6604 17255
rect 6552 17212 6604 17221
rect 2228 17076 2280 17128
rect 3516 17144 3568 17196
rect 6644 17144 6696 17196
rect 7932 17212 7984 17264
rect 8576 17212 8628 17264
rect 9864 17255 9916 17264
rect 9864 17221 9873 17255
rect 9873 17221 9907 17255
rect 9907 17221 9916 17255
rect 9864 17212 9916 17221
rect 10876 17212 10928 17264
rect 9588 17187 9640 17196
rect 9588 17153 9597 17187
rect 9597 17153 9631 17187
rect 9631 17153 9640 17187
rect 9588 17144 9640 17153
rect 11428 17144 11480 17196
rect 11704 17187 11756 17196
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 3884 17119 3936 17128
rect 3884 17085 3893 17119
rect 3893 17085 3927 17119
rect 3927 17085 3936 17119
rect 3884 17076 3936 17085
rect 11336 17119 11388 17128
rect 11336 17085 11345 17119
rect 11345 17085 11379 17119
rect 11379 17085 11388 17119
rect 11336 17076 11388 17085
rect 3516 17008 3568 17060
rect 10968 17008 11020 17060
rect 12256 17187 12308 17196
rect 12256 17153 12265 17187
rect 12265 17153 12299 17187
rect 12299 17153 12308 17187
rect 14924 17212 14976 17264
rect 12256 17144 12308 17153
rect 13728 17144 13780 17196
rect 15200 17187 15252 17196
rect 15200 17153 15210 17187
rect 15210 17153 15244 17187
rect 15244 17153 15252 17187
rect 15200 17144 15252 17153
rect 17132 17144 17184 17196
rect 17592 17187 17644 17196
rect 17592 17153 17601 17187
rect 17601 17153 17635 17187
rect 17635 17153 17644 17187
rect 17592 17144 17644 17153
rect 12440 17076 12492 17128
rect 17776 17144 17828 17196
rect 18144 17187 18196 17196
rect 18696 17212 18748 17264
rect 18144 17153 18183 17187
rect 18183 17153 18196 17187
rect 18144 17144 18196 17153
rect 17868 17008 17920 17060
rect 1400 16983 1452 16992
rect 1400 16949 1409 16983
rect 1409 16949 1443 16983
rect 1443 16949 1452 16983
rect 1400 16940 1452 16949
rect 2044 16983 2096 16992
rect 2044 16949 2053 16983
rect 2053 16949 2087 16983
rect 2087 16949 2096 16983
rect 2044 16940 2096 16949
rect 2780 16940 2832 16992
rect 3792 16940 3844 16992
rect 6092 16983 6144 16992
rect 6092 16949 6101 16983
rect 6101 16949 6135 16983
rect 6135 16949 6144 16983
rect 6092 16940 6144 16949
rect 17316 16940 17368 16992
rect 18420 16940 18472 16992
rect 2350 16838 2402 16890
rect 2414 16838 2466 16890
rect 2478 16838 2530 16890
rect 2542 16838 2594 16890
rect 2606 16838 2658 16890
rect 1584 16736 1636 16788
rect 1676 16736 1728 16788
rect 3884 16668 3936 16720
rect 1676 16643 1728 16652
rect 1676 16609 1685 16643
rect 1685 16609 1719 16643
rect 1719 16609 1728 16643
rect 1676 16600 1728 16609
rect 2044 16600 2096 16652
rect 3792 16600 3844 16652
rect 6460 16779 6512 16788
rect 6460 16745 6469 16779
rect 6469 16745 6503 16779
rect 6503 16745 6512 16779
rect 6460 16736 6512 16745
rect 1584 16575 1636 16584
rect 1584 16541 1593 16575
rect 1593 16541 1627 16575
rect 1627 16541 1636 16575
rect 1584 16532 1636 16541
rect 5724 16600 5776 16652
rect 6552 16643 6604 16652
rect 6552 16609 6561 16643
rect 6561 16609 6595 16643
rect 6595 16609 6604 16643
rect 6552 16600 6604 16609
rect 9588 16600 9640 16652
rect 12624 16736 12676 16788
rect 12716 16736 12768 16788
rect 13728 16736 13780 16788
rect 10968 16643 11020 16652
rect 10968 16609 10977 16643
rect 10977 16609 11011 16643
rect 11011 16609 11020 16643
rect 10968 16600 11020 16609
rect 11428 16600 11480 16652
rect 2780 16396 2832 16448
rect 4620 16575 4672 16584
rect 4620 16541 4629 16575
rect 4629 16541 4663 16575
rect 4663 16541 4672 16575
rect 4620 16532 4672 16541
rect 6092 16532 6144 16584
rect 6368 16532 6420 16584
rect 4896 16464 4948 16516
rect 8300 16507 8352 16516
rect 8300 16473 8309 16507
rect 8309 16473 8343 16507
rect 8343 16473 8352 16507
rect 8300 16464 8352 16473
rect 9220 16532 9272 16584
rect 12716 16575 12768 16584
rect 12716 16541 12725 16575
rect 12725 16541 12759 16575
rect 12759 16541 12768 16575
rect 12716 16532 12768 16541
rect 18696 16736 18748 16788
rect 15844 16600 15896 16652
rect 17316 16643 17368 16652
rect 17316 16609 17325 16643
rect 17325 16609 17359 16643
rect 17359 16609 17368 16643
rect 17316 16600 17368 16609
rect 3424 16439 3476 16448
rect 3424 16405 3433 16439
rect 3433 16405 3467 16439
rect 3467 16405 3476 16439
rect 3424 16396 3476 16405
rect 4068 16439 4120 16448
rect 4068 16405 4077 16439
rect 4077 16405 4111 16439
rect 4111 16405 4120 16439
rect 4068 16396 4120 16405
rect 4620 16396 4672 16448
rect 6368 16396 6420 16448
rect 6644 16396 6696 16448
rect 8668 16396 8720 16448
rect 9496 16396 9548 16448
rect 14924 16575 14976 16584
rect 14924 16541 14933 16575
rect 14933 16541 14967 16575
rect 14967 16541 14976 16575
rect 14924 16532 14976 16541
rect 15016 16575 15068 16584
rect 15016 16541 15026 16575
rect 15026 16541 15060 16575
rect 15060 16541 15068 16575
rect 15016 16532 15068 16541
rect 18420 16532 18472 16584
rect 12256 16396 12308 16448
rect 12440 16439 12492 16448
rect 12440 16405 12449 16439
rect 12449 16405 12483 16439
rect 12483 16405 12492 16439
rect 12440 16396 12492 16405
rect 14464 16396 14516 16448
rect 14556 16439 14608 16448
rect 14556 16405 14565 16439
rect 14565 16405 14599 16439
rect 14599 16405 14608 16439
rect 14556 16396 14608 16405
rect 16212 16396 16264 16448
rect 17132 16396 17184 16448
rect 3010 16294 3062 16346
rect 3074 16294 3126 16346
rect 3138 16294 3190 16346
rect 3202 16294 3254 16346
rect 3266 16294 3318 16346
rect 2228 16192 2280 16244
rect 2780 16235 2832 16244
rect 2780 16201 2789 16235
rect 2789 16201 2823 16235
rect 2823 16201 2832 16235
rect 2780 16192 2832 16201
rect 4896 16235 4948 16244
rect 4896 16201 4905 16235
rect 4905 16201 4939 16235
rect 4939 16201 4948 16235
rect 4896 16192 4948 16201
rect 1584 16124 1636 16176
rect 848 16056 900 16108
rect 3424 16124 3476 16176
rect 4068 16124 4120 16176
rect 8392 16192 8444 16244
rect 9220 16235 9272 16244
rect 9220 16201 9229 16235
rect 9229 16201 9263 16235
rect 9263 16201 9272 16235
rect 9220 16192 9272 16201
rect 12624 16192 12676 16244
rect 15844 16192 15896 16244
rect 18512 16192 18564 16244
rect 2136 16099 2188 16108
rect 2136 16065 2146 16099
rect 2146 16065 2180 16099
rect 2180 16065 2188 16099
rect 2136 16056 2188 16065
rect 2688 16099 2740 16108
rect 2688 16065 2697 16099
rect 2697 16065 2731 16099
rect 2731 16065 2740 16099
rect 2688 16056 2740 16065
rect 2872 16056 2924 16108
rect 6920 16056 6972 16108
rect 8484 16124 8536 16176
rect 13268 16124 13320 16176
rect 17500 16124 17552 16176
rect 7380 16099 7432 16108
rect 7380 16065 7389 16099
rect 7389 16065 7423 16099
rect 7423 16065 7432 16099
rect 7380 16056 7432 16065
rect 9496 16099 9548 16108
rect 9496 16065 9505 16099
rect 9505 16065 9539 16099
rect 9539 16065 9548 16099
rect 9496 16056 9548 16065
rect 14188 16099 14240 16108
rect 14188 16065 14197 16099
rect 14197 16065 14231 16099
rect 14231 16065 14240 16099
rect 14188 16056 14240 16065
rect 15936 16056 15988 16108
rect 18788 16099 18840 16108
rect 18788 16065 18797 16099
rect 18797 16065 18831 16099
rect 18831 16065 18840 16099
rect 18788 16056 18840 16065
rect 6552 15988 6604 16040
rect 8116 15988 8168 16040
rect 9680 15963 9732 15972
rect 9680 15929 9689 15963
rect 9689 15929 9723 15963
rect 9723 15929 9732 15963
rect 9680 15920 9732 15929
rect 1768 15852 1820 15904
rect 2688 15852 2740 15904
rect 5816 15852 5868 15904
rect 7288 15895 7340 15904
rect 7288 15861 7297 15895
rect 7297 15861 7331 15895
rect 7331 15861 7340 15895
rect 7288 15852 7340 15861
rect 14096 15988 14148 16040
rect 17316 15988 17368 16040
rect 13360 15852 13412 15904
rect 14372 15852 14424 15904
rect 18144 15852 18196 15904
rect 2350 15750 2402 15802
rect 2414 15750 2466 15802
rect 2478 15750 2530 15802
rect 2542 15750 2594 15802
rect 2606 15750 2658 15802
rect 3424 15444 3476 15496
rect 5816 15487 5868 15496
rect 5816 15453 5825 15487
rect 5825 15453 5859 15487
rect 5859 15453 5868 15487
rect 6644 15648 6696 15700
rect 8116 15648 8168 15700
rect 8484 15648 8536 15700
rect 11520 15648 11572 15700
rect 13268 15648 13320 15700
rect 15016 15648 15068 15700
rect 17132 15691 17184 15700
rect 17132 15657 17141 15691
rect 17141 15657 17175 15691
rect 17175 15657 17184 15691
rect 17132 15648 17184 15657
rect 17500 15691 17552 15700
rect 17500 15657 17509 15691
rect 17509 15657 17543 15691
rect 17543 15657 17552 15691
rect 17500 15648 17552 15657
rect 6552 15512 6604 15564
rect 5816 15444 5868 15453
rect 12716 15512 12768 15564
rect 1400 15351 1452 15360
rect 1400 15317 1409 15351
rect 1409 15317 1443 15351
rect 1443 15317 1452 15351
rect 1400 15308 1452 15317
rect 2136 15308 2188 15360
rect 2688 15308 2740 15360
rect 5724 15351 5776 15360
rect 5724 15317 5733 15351
rect 5733 15317 5767 15351
rect 5767 15317 5776 15351
rect 5724 15308 5776 15317
rect 7196 15308 7248 15360
rect 9312 15419 9364 15428
rect 9312 15385 9321 15419
rect 9321 15385 9355 15419
rect 9355 15385 9364 15419
rect 9312 15376 9364 15385
rect 8668 15308 8720 15360
rect 12624 15444 12676 15496
rect 17592 15580 17644 15632
rect 15936 15555 15988 15564
rect 15936 15521 15945 15555
rect 15945 15521 15979 15555
rect 15979 15521 15988 15555
rect 15936 15512 15988 15521
rect 16212 15555 16264 15564
rect 16212 15521 16221 15555
rect 16221 15521 16255 15555
rect 16255 15521 16264 15555
rect 16212 15512 16264 15521
rect 13728 15444 13780 15496
rect 14556 15444 14608 15496
rect 14372 15308 14424 15360
rect 16764 15487 16816 15496
rect 16764 15453 16773 15487
rect 16773 15453 16807 15487
rect 16807 15453 16816 15487
rect 16764 15444 16816 15453
rect 17500 15444 17552 15496
rect 17868 15444 17920 15496
rect 18328 15444 18380 15496
rect 18512 15376 18564 15428
rect 17316 15351 17368 15360
rect 17316 15317 17325 15351
rect 17325 15317 17359 15351
rect 17359 15317 17368 15351
rect 17316 15308 17368 15317
rect 18788 15351 18840 15360
rect 18788 15317 18797 15351
rect 18797 15317 18831 15351
rect 18831 15317 18840 15351
rect 18788 15308 18840 15317
rect 3010 15206 3062 15258
rect 3074 15206 3126 15258
rect 3138 15206 3190 15258
rect 3202 15206 3254 15258
rect 3266 15206 3318 15258
rect 1860 15104 1912 15156
rect 3424 15104 3476 15156
rect 2964 15036 3016 15088
rect 5724 15036 5776 15088
rect 7012 15036 7064 15088
rect 7196 15147 7248 15156
rect 7196 15113 7205 15147
rect 7205 15113 7239 15147
rect 7239 15113 7248 15147
rect 7196 15104 7248 15113
rect 7288 15104 7340 15156
rect 14096 15147 14148 15156
rect 14096 15113 14105 15147
rect 14105 15113 14139 15147
rect 14139 15113 14148 15147
rect 14096 15104 14148 15113
rect 14464 15147 14516 15156
rect 14464 15113 14473 15147
rect 14473 15113 14507 15147
rect 14507 15113 14516 15147
rect 14464 15104 14516 15113
rect 2780 14968 2832 15020
rect 1676 14943 1728 14952
rect 1676 14909 1685 14943
rect 1685 14909 1719 14943
rect 1719 14909 1728 14943
rect 1676 14900 1728 14909
rect 1768 14900 1820 14952
rect 2688 14900 2740 14952
rect 3700 15011 3752 15020
rect 3700 14977 3709 15011
rect 3709 14977 3743 15011
rect 3743 14977 3752 15011
rect 3700 14968 3752 14977
rect 3792 15011 3844 15020
rect 3792 14977 3801 15011
rect 3801 14977 3835 15011
rect 3835 14977 3844 15011
rect 3792 14968 3844 14977
rect 5632 15011 5684 15020
rect 5632 14977 5641 15011
rect 5641 14977 5675 15011
rect 5675 14977 5684 15011
rect 5632 14968 5684 14977
rect 9312 15036 9364 15088
rect 11428 15036 11480 15088
rect 8116 14968 8168 15020
rect 11796 15011 11848 15020
rect 11796 14977 11805 15011
rect 11805 14977 11839 15011
rect 11839 14977 11848 15011
rect 11796 14968 11848 14977
rect 17316 15036 17368 15088
rect 14372 14968 14424 15020
rect 17040 14968 17092 15020
rect 4068 14943 4120 14952
rect 4068 14909 4077 14943
rect 4077 14909 4111 14943
rect 4111 14909 4120 14943
rect 4068 14900 4120 14909
rect 4528 14900 4580 14952
rect 15476 14943 15528 14952
rect 15476 14909 15485 14943
rect 15485 14909 15519 14943
rect 15519 14909 15528 14943
rect 15476 14900 15528 14909
rect 15660 14943 15712 14952
rect 15660 14909 15669 14943
rect 15669 14909 15703 14943
rect 15703 14909 15712 14943
rect 15660 14900 15712 14909
rect 17776 15011 17828 15020
rect 17776 14977 17785 15011
rect 17785 14977 17819 15011
rect 17819 14977 17828 15011
rect 17776 14968 17828 14977
rect 18144 15011 18196 15020
rect 18144 14977 18152 15011
rect 18152 14977 18186 15011
rect 18186 14977 18196 15011
rect 18144 14968 18196 14977
rect 18236 15011 18288 15020
rect 18236 14977 18245 15011
rect 18245 14977 18279 15011
rect 18279 14977 18288 15011
rect 18236 14968 18288 14977
rect 18880 14968 18932 15020
rect 17960 14832 18012 14884
rect 3608 14807 3660 14816
rect 3608 14773 3617 14807
rect 3617 14773 3651 14807
rect 3651 14773 3660 14807
rect 3608 14764 3660 14773
rect 5540 14807 5592 14816
rect 5540 14773 5549 14807
rect 5549 14773 5583 14807
rect 5583 14773 5592 14807
rect 5540 14764 5592 14773
rect 6920 14807 6972 14816
rect 6920 14773 6929 14807
rect 6929 14773 6963 14807
rect 6963 14773 6972 14807
rect 6920 14764 6972 14773
rect 17316 14764 17368 14816
rect 17408 14764 17460 14816
rect 2350 14662 2402 14714
rect 2414 14662 2466 14714
rect 2478 14662 2530 14714
rect 2542 14662 2594 14714
rect 2606 14662 2658 14714
rect 2780 14560 2832 14612
rect 4068 14560 4120 14612
rect 14648 14560 14700 14612
rect 1952 14492 2004 14544
rect 3516 14492 3568 14544
rect 3700 14492 3752 14544
rect 13360 14492 13412 14544
rect 1676 14424 1728 14476
rect 1768 14399 1820 14408
rect 1768 14365 1777 14399
rect 1777 14365 1811 14399
rect 1811 14365 1820 14399
rect 1768 14356 1820 14365
rect 2136 14356 2188 14408
rect 3792 14424 3844 14476
rect 5632 14424 5684 14476
rect 11428 14424 11480 14476
rect 3608 14288 3660 14340
rect 4344 14399 4396 14408
rect 4344 14365 4353 14399
rect 4353 14365 4387 14399
rect 4387 14365 4396 14399
rect 4344 14356 4396 14365
rect 4528 14399 4580 14408
rect 4528 14365 4537 14399
rect 4537 14365 4571 14399
rect 4571 14365 4580 14399
rect 4528 14356 4580 14365
rect 8300 14356 8352 14408
rect 10968 14356 11020 14408
rect 13728 14356 13780 14408
rect 14372 14356 14424 14408
rect 16948 14424 17000 14476
rect 17316 14467 17368 14476
rect 17316 14433 17325 14467
rect 17325 14433 17359 14467
rect 17359 14433 17368 14467
rect 17316 14424 17368 14433
rect 5540 14288 5592 14340
rect 14648 14399 14700 14408
rect 14648 14365 14657 14399
rect 14657 14365 14691 14399
rect 14691 14365 14700 14399
rect 14648 14356 14700 14365
rect 16856 14356 16908 14408
rect 16028 14288 16080 14340
rect 18052 14288 18104 14340
rect 1676 14263 1728 14272
rect 1676 14229 1685 14263
rect 1685 14229 1719 14263
rect 1719 14229 1728 14263
rect 1676 14220 1728 14229
rect 1768 14220 1820 14272
rect 3516 14220 3568 14272
rect 4528 14220 4580 14272
rect 14280 14220 14332 14272
rect 14464 14263 14516 14272
rect 14464 14229 14473 14263
rect 14473 14229 14507 14263
rect 14507 14229 14516 14263
rect 14464 14220 14516 14229
rect 15384 14220 15436 14272
rect 16488 14263 16540 14272
rect 16488 14229 16497 14263
rect 16497 14229 16531 14263
rect 16531 14229 16540 14263
rect 16488 14220 16540 14229
rect 18236 14220 18288 14272
rect 3010 14118 3062 14170
rect 3074 14118 3126 14170
rect 3138 14118 3190 14170
rect 3202 14118 3254 14170
rect 3266 14118 3318 14170
rect 1676 14016 1728 14068
rect 17408 14016 17460 14068
rect 18052 14059 18104 14068
rect 18052 14025 18061 14059
rect 18061 14025 18095 14059
rect 18095 14025 18104 14059
rect 18052 14016 18104 14025
rect 18788 14059 18840 14068
rect 18788 14025 18797 14059
rect 18797 14025 18831 14059
rect 18831 14025 18840 14059
rect 18788 14016 18840 14025
rect 1032 13948 1084 14000
rect 1492 13923 1544 13932
rect 1492 13889 1501 13923
rect 1501 13889 1535 13923
rect 1535 13889 1544 13923
rect 1492 13880 1544 13889
rect 2688 13948 2740 14000
rect 2136 13880 2188 13932
rect 3884 13880 3936 13932
rect 4252 13880 4304 13932
rect 4068 13812 4120 13864
rect 4620 13880 4672 13932
rect 13360 13923 13412 13932
rect 13360 13889 13369 13923
rect 13369 13889 13403 13923
rect 13403 13889 13412 13923
rect 13360 13880 13412 13889
rect 16580 13880 16632 13932
rect 16764 13880 16816 13932
rect 1768 13744 1820 13796
rect 5540 13855 5592 13864
rect 5540 13821 5549 13855
rect 5549 13821 5583 13855
rect 5583 13821 5592 13855
rect 5540 13812 5592 13821
rect 5816 13855 5868 13864
rect 5816 13821 5825 13855
rect 5825 13821 5859 13855
rect 5859 13821 5868 13855
rect 5816 13812 5868 13821
rect 14372 13812 14424 13864
rect 16120 13812 16172 13864
rect 17500 13812 17552 13864
rect 18420 13880 18472 13932
rect 18604 13923 18656 13932
rect 18604 13889 18613 13923
rect 18613 13889 18647 13923
rect 18647 13889 18656 13923
rect 18604 13880 18656 13889
rect 6000 13744 6052 13796
rect 3148 13676 3200 13728
rect 4620 13676 4672 13728
rect 17040 13719 17092 13728
rect 17040 13685 17049 13719
rect 17049 13685 17083 13719
rect 17083 13685 17092 13719
rect 17040 13676 17092 13685
rect 17224 13719 17276 13728
rect 17224 13685 17233 13719
rect 17233 13685 17267 13719
rect 17267 13685 17276 13719
rect 17224 13676 17276 13685
rect 2350 13574 2402 13626
rect 2414 13574 2466 13626
rect 2478 13574 2530 13626
rect 2542 13574 2594 13626
rect 2606 13574 2658 13626
rect 3792 13515 3844 13524
rect 3792 13481 3801 13515
rect 3801 13481 3835 13515
rect 3835 13481 3844 13515
rect 3792 13472 3844 13481
rect 5816 13472 5868 13524
rect 6000 13472 6052 13524
rect 13912 13472 13964 13524
rect 15108 13472 15160 13524
rect 16028 13515 16080 13524
rect 16028 13481 16037 13515
rect 16037 13481 16071 13515
rect 16071 13481 16080 13515
rect 16028 13472 16080 13481
rect 18604 13515 18656 13524
rect 18604 13481 18613 13515
rect 18613 13481 18647 13515
rect 18647 13481 18656 13515
rect 18604 13472 18656 13481
rect 1860 13379 1912 13388
rect 1860 13345 1869 13379
rect 1869 13345 1903 13379
rect 1903 13345 1912 13379
rect 1860 13336 1912 13345
rect 4620 13379 4672 13388
rect 4620 13345 4629 13379
rect 4629 13345 4663 13379
rect 4663 13345 4672 13379
rect 4620 13336 4672 13345
rect 1584 13175 1636 13184
rect 1584 13141 1593 13175
rect 1593 13141 1627 13175
rect 1627 13141 1636 13175
rect 1584 13132 1636 13141
rect 4068 13311 4120 13320
rect 4068 13277 4077 13311
rect 4077 13277 4111 13311
rect 4111 13277 4120 13311
rect 4068 13268 4120 13277
rect 2136 13243 2188 13252
rect 2136 13209 2145 13243
rect 2145 13209 2179 13243
rect 2179 13209 2188 13243
rect 2136 13200 2188 13209
rect 3148 13200 3200 13252
rect 3884 13200 3936 13252
rect 6368 13311 6420 13320
rect 6368 13277 6377 13311
rect 6377 13277 6411 13311
rect 6411 13277 6420 13311
rect 6368 13268 6420 13277
rect 6644 13268 6696 13320
rect 14464 13336 14516 13388
rect 17224 13336 17276 13388
rect 14004 13268 14056 13320
rect 10968 13200 11020 13252
rect 14188 13268 14240 13320
rect 15752 13268 15804 13320
rect 16120 13311 16172 13320
rect 16120 13277 16129 13311
rect 16129 13277 16163 13311
rect 16163 13277 16172 13311
rect 16120 13268 16172 13277
rect 15108 13200 15160 13252
rect 16856 13200 16908 13252
rect 2872 13132 2924 13184
rect 3976 13175 4028 13184
rect 3976 13141 3985 13175
rect 3985 13141 4019 13175
rect 4019 13141 4028 13175
rect 3976 13132 4028 13141
rect 13176 13132 13228 13184
rect 18420 13132 18472 13184
rect 3010 13030 3062 13082
rect 3074 13030 3126 13082
rect 3138 13030 3190 13082
rect 3202 13030 3254 13082
rect 3266 13030 3318 13082
rect 1216 12928 1268 12980
rect 2136 12928 2188 12980
rect 13360 12928 13412 12980
rect 13912 12928 13964 12980
rect 14004 12928 14056 12980
rect 15476 12928 15528 12980
rect 15660 12971 15712 12980
rect 15660 12937 15669 12971
rect 15669 12937 15703 12971
rect 15703 12937 15712 12971
rect 15660 12928 15712 12937
rect 18328 12971 18380 12980
rect 18328 12937 18337 12971
rect 18337 12937 18371 12971
rect 18371 12937 18380 12971
rect 18328 12928 18380 12937
rect 18512 12928 18564 12980
rect 1584 12835 1636 12844
rect 1584 12801 1593 12835
rect 1593 12801 1627 12835
rect 1627 12801 1636 12835
rect 1584 12792 1636 12801
rect 1676 12835 1728 12844
rect 1676 12801 1685 12835
rect 1685 12801 1719 12835
rect 1719 12801 1728 12835
rect 1676 12792 1728 12801
rect 1768 12792 1820 12844
rect 2872 12835 2924 12844
rect 2872 12801 2881 12835
rect 2881 12801 2915 12835
rect 2915 12801 2924 12835
rect 2872 12792 2924 12801
rect 3424 12860 3476 12912
rect 5356 12860 5408 12912
rect 3976 12792 4028 12844
rect 14280 12792 14332 12844
rect 15200 12792 15252 12844
rect 16488 12792 16540 12844
rect 18144 12835 18196 12844
rect 18144 12801 18153 12835
rect 18153 12801 18187 12835
rect 18187 12801 18196 12835
rect 18144 12792 18196 12801
rect 18788 12835 18840 12844
rect 18788 12801 18797 12835
rect 18797 12801 18831 12835
rect 18831 12801 18840 12835
rect 18788 12792 18840 12801
rect 4068 12724 4120 12776
rect 13176 12767 13228 12776
rect 13176 12733 13185 12767
rect 13185 12733 13219 12767
rect 13219 12733 13228 12767
rect 13176 12724 13228 12733
rect 7012 12588 7064 12640
rect 2350 12486 2402 12538
rect 2414 12486 2466 12538
rect 2478 12486 2530 12538
rect 2542 12486 2594 12538
rect 2606 12486 2658 12538
rect 11888 12384 11940 12436
rect 15108 12384 15160 12436
rect 13912 12291 13964 12300
rect 13912 12257 13921 12291
rect 13921 12257 13955 12291
rect 13955 12257 13964 12291
rect 13912 12248 13964 12257
rect 11888 12155 11940 12164
rect 11888 12121 11897 12155
rect 11897 12121 11931 12155
rect 11931 12121 11940 12155
rect 11888 12112 11940 12121
rect 12992 12112 13044 12164
rect 3884 12044 3936 12096
rect 4436 12044 4488 12096
rect 14372 12155 14424 12164
rect 14372 12121 14381 12155
rect 14381 12121 14415 12155
rect 14415 12121 14424 12155
rect 14372 12112 14424 12121
rect 15108 12112 15160 12164
rect 17408 12112 17460 12164
rect 18144 12223 18196 12232
rect 18144 12189 18153 12223
rect 18153 12189 18187 12223
rect 18187 12189 18196 12223
rect 18144 12180 18196 12189
rect 18696 12180 18748 12232
rect 18788 12223 18840 12232
rect 18788 12189 18797 12223
rect 18797 12189 18831 12223
rect 18831 12189 18840 12223
rect 18788 12180 18840 12189
rect 15384 12044 15436 12096
rect 15660 12044 15712 12096
rect 17592 12044 17644 12096
rect 3010 11942 3062 11994
rect 3074 11942 3126 11994
rect 3138 11942 3190 11994
rect 3202 11942 3254 11994
rect 3266 11942 3318 11994
rect 1768 11772 1820 11824
rect 2136 11772 2188 11824
rect 4160 11840 4212 11892
rect 4804 11840 4856 11892
rect 12992 11883 13044 11892
rect 12992 11849 13001 11883
rect 13001 11849 13035 11883
rect 13035 11849 13044 11883
rect 12992 11840 13044 11849
rect 15108 11883 15160 11892
rect 15108 11849 15117 11883
rect 15117 11849 15151 11883
rect 15151 11849 15160 11883
rect 15108 11840 15160 11849
rect 18696 11883 18748 11892
rect 18696 11849 18705 11883
rect 18705 11849 18739 11883
rect 18739 11849 18748 11883
rect 18696 11840 18748 11849
rect 3884 11704 3936 11756
rect 4068 11747 4120 11756
rect 4068 11713 4077 11747
rect 4077 11713 4111 11747
rect 4111 11713 4120 11747
rect 4068 11704 4120 11713
rect 4160 11747 4212 11756
rect 4160 11713 4169 11747
rect 4169 11713 4203 11747
rect 4203 11713 4212 11747
rect 4160 11704 4212 11713
rect 5080 11772 5132 11824
rect 17500 11772 17552 11824
rect 17960 11772 18012 11824
rect 4436 11747 4488 11756
rect 4436 11713 4445 11747
rect 4445 11713 4479 11747
rect 4479 11713 4488 11747
rect 4436 11704 4488 11713
rect 4804 11747 4856 11756
rect 4804 11713 4813 11747
rect 4813 11713 4847 11747
rect 4847 11713 4856 11747
rect 4804 11704 4856 11713
rect 4988 11747 5040 11756
rect 4988 11713 4997 11747
rect 4997 11713 5031 11747
rect 5031 11713 5040 11747
rect 4988 11704 5040 11713
rect 6368 11704 6420 11756
rect 1768 11636 1820 11688
rect 3148 11543 3200 11552
rect 3148 11509 3157 11543
rect 3157 11509 3191 11543
rect 3191 11509 3200 11543
rect 3148 11500 3200 11509
rect 4160 11500 4212 11552
rect 4712 11679 4764 11688
rect 4712 11645 4721 11679
rect 4721 11645 4755 11679
rect 4755 11645 4764 11679
rect 4712 11636 4764 11645
rect 4896 11543 4948 11552
rect 4896 11509 4905 11543
rect 4905 11509 4939 11543
rect 4939 11509 4948 11543
rect 4896 11500 4948 11509
rect 5080 11543 5132 11552
rect 5080 11509 5089 11543
rect 5089 11509 5123 11543
rect 5123 11509 5132 11543
rect 5080 11500 5132 11509
rect 5264 11500 5316 11552
rect 10600 11543 10652 11552
rect 10600 11509 10609 11543
rect 10609 11509 10643 11543
rect 10643 11509 10652 11543
rect 10600 11500 10652 11509
rect 10968 11500 11020 11552
rect 15200 11704 15252 11756
rect 15660 11704 15712 11756
rect 16948 11747 17000 11756
rect 16948 11713 16957 11747
rect 16957 11713 16991 11747
rect 16991 11713 17000 11747
rect 16948 11704 17000 11713
rect 15844 11679 15896 11688
rect 15844 11645 15853 11679
rect 15853 11645 15887 11679
rect 15887 11645 15896 11679
rect 15844 11636 15896 11645
rect 17224 11679 17276 11688
rect 17224 11645 17233 11679
rect 17233 11645 17267 11679
rect 17267 11645 17276 11679
rect 17224 11636 17276 11645
rect 15936 11568 15988 11620
rect 15752 11500 15804 11552
rect 2350 11398 2402 11450
rect 2414 11398 2466 11450
rect 2478 11398 2530 11450
rect 2542 11398 2594 11450
rect 2606 11398 2658 11450
rect 2136 11339 2188 11348
rect 2136 11305 2145 11339
rect 2145 11305 2179 11339
rect 2179 11305 2188 11339
rect 2136 11296 2188 11305
rect 4068 11296 4120 11348
rect 4712 11296 4764 11348
rect 3148 11271 3200 11280
rect 3148 11237 3157 11271
rect 3157 11237 3191 11271
rect 3191 11237 3200 11271
rect 3148 11228 3200 11237
rect 3792 11228 3844 11280
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 2228 11135 2280 11144
rect 2228 11101 2237 11135
rect 2237 11101 2271 11135
rect 2271 11101 2280 11135
rect 2228 11092 2280 11101
rect 2780 11067 2832 11076
rect 2780 11033 2789 11067
rect 2789 11033 2823 11067
rect 2823 11033 2832 11067
rect 2780 11024 2832 11033
rect 3516 11024 3568 11076
rect 1584 10999 1636 11008
rect 1584 10965 1593 10999
rect 1593 10965 1627 10999
rect 1627 10965 1636 10999
rect 1584 10956 1636 10965
rect 3884 11135 3936 11144
rect 3884 11101 3893 11135
rect 3893 11101 3927 11135
rect 3927 11101 3936 11135
rect 3884 11092 3936 11101
rect 4804 11228 4856 11280
rect 4896 11228 4948 11280
rect 5356 11296 5408 11348
rect 5540 11296 5592 11348
rect 6368 11296 6420 11348
rect 5816 11160 5868 11212
rect 6828 11160 6880 11212
rect 4252 11092 4304 11144
rect 4896 11135 4948 11144
rect 4896 11101 4905 11135
rect 4905 11101 4939 11135
rect 4939 11101 4948 11135
rect 4896 11092 4948 11101
rect 5080 11092 5132 11144
rect 14372 11092 14424 11144
rect 15384 11228 15436 11280
rect 16488 11228 16540 11280
rect 17224 11296 17276 11348
rect 17960 11296 18012 11348
rect 17408 11228 17460 11280
rect 15568 11092 15620 11144
rect 15752 11135 15804 11144
rect 15752 11101 15761 11135
rect 15761 11101 15795 11135
rect 15795 11101 15804 11135
rect 15752 11092 15804 11101
rect 17408 11135 17460 11144
rect 17408 11101 17417 11135
rect 17417 11101 17451 11135
rect 17451 11101 17460 11135
rect 17408 11092 17460 11101
rect 17500 11135 17552 11144
rect 17500 11101 17509 11135
rect 17509 11101 17543 11135
rect 17543 11101 17552 11135
rect 17500 11092 17552 11101
rect 17592 11135 17644 11144
rect 17592 11101 17601 11135
rect 17601 11101 17635 11135
rect 17635 11101 17644 11135
rect 17592 11092 17644 11101
rect 17776 11135 17828 11144
rect 17776 11101 17785 11135
rect 17785 11101 17819 11135
rect 17819 11101 17828 11135
rect 17776 11092 17828 11101
rect 18420 11092 18472 11144
rect 18788 11135 18840 11144
rect 18788 11101 18797 11135
rect 18797 11101 18831 11135
rect 18831 11101 18840 11135
rect 18788 11092 18840 11101
rect 6092 11024 6144 11076
rect 15660 11067 15712 11076
rect 15660 11033 15669 11067
rect 15669 11033 15703 11067
rect 15703 11033 15712 11067
rect 15660 11024 15712 11033
rect 6828 10956 6880 11008
rect 15476 10999 15528 11008
rect 15476 10965 15485 10999
rect 15485 10965 15519 10999
rect 15519 10965 15528 10999
rect 15476 10956 15528 10965
rect 16856 10956 16908 11008
rect 3010 10854 3062 10906
rect 3074 10854 3126 10906
rect 3138 10854 3190 10906
rect 3202 10854 3254 10906
rect 3266 10854 3318 10906
rect 3884 10752 3936 10804
rect 4528 10752 4580 10804
rect 4896 10752 4948 10804
rect 1584 10684 1636 10736
rect 2228 10684 2280 10736
rect 5264 10684 5316 10736
rect 5540 10727 5592 10736
rect 5540 10693 5549 10727
rect 5549 10693 5583 10727
rect 5583 10693 5592 10727
rect 5540 10684 5592 10693
rect 6092 10752 6144 10804
rect 6828 10795 6880 10804
rect 6828 10761 6837 10795
rect 6837 10761 6871 10795
rect 6871 10761 6880 10795
rect 6828 10752 6880 10761
rect 15844 10752 15896 10804
rect 5816 10659 5868 10668
rect 5816 10625 5825 10659
rect 5825 10625 5859 10659
rect 5859 10625 5868 10659
rect 5816 10616 5868 10625
rect 15660 10616 15712 10668
rect 18328 10616 18380 10668
rect 1400 10591 1452 10600
rect 1400 10557 1409 10591
rect 1409 10557 1443 10591
rect 1443 10557 1452 10591
rect 1400 10548 1452 10557
rect 4988 10548 5040 10600
rect 6736 10548 6788 10600
rect 14188 10548 14240 10600
rect 15200 10548 15252 10600
rect 17960 10548 18012 10600
rect 18604 10412 18656 10464
rect 18788 10455 18840 10464
rect 18788 10421 18797 10455
rect 18797 10421 18831 10455
rect 18831 10421 18840 10455
rect 18788 10412 18840 10421
rect 2350 10310 2402 10362
rect 2414 10310 2466 10362
rect 2478 10310 2530 10362
rect 2542 10310 2594 10362
rect 2606 10310 2658 10362
rect 2228 10208 2280 10260
rect 15200 10251 15252 10260
rect 15200 10217 15209 10251
rect 15209 10217 15243 10251
rect 15243 10217 15252 10251
rect 15200 10208 15252 10217
rect 18328 10251 18380 10260
rect 18328 10217 18337 10251
rect 18337 10217 18371 10251
rect 18371 10217 18380 10251
rect 18328 10208 18380 10217
rect 848 10072 900 10124
rect 8208 10072 8260 10124
rect 16856 10115 16908 10124
rect 16856 10081 16865 10115
rect 16865 10081 16899 10115
rect 16899 10081 16908 10115
rect 16856 10072 16908 10081
rect 2136 10004 2188 10056
rect 15476 10004 15528 10056
rect 15844 10004 15896 10056
rect 16580 10047 16632 10056
rect 16580 10013 16589 10047
rect 16589 10013 16623 10047
rect 16623 10013 16632 10047
rect 16580 10004 16632 10013
rect 18420 10047 18472 10056
rect 18420 10013 18429 10047
rect 18429 10013 18463 10047
rect 18463 10013 18472 10047
rect 18420 10004 18472 10013
rect 16856 9936 16908 9988
rect 3010 9766 3062 9818
rect 3074 9766 3126 9818
rect 3138 9766 3190 9818
rect 3202 9766 3254 9818
rect 3266 9766 3318 9818
rect 2872 9596 2924 9648
rect 4160 9639 4212 9648
rect 4160 9605 4169 9639
rect 4169 9605 4203 9639
rect 4203 9605 4212 9639
rect 4160 9596 4212 9605
rect 8116 9596 8168 9648
rect 10600 9596 10652 9648
rect 12532 9596 12584 9648
rect 17408 9596 17460 9648
rect 848 9528 900 9580
rect 1492 9528 1544 9580
rect 5908 9571 5960 9580
rect 5908 9537 5917 9571
rect 5917 9537 5951 9571
rect 5951 9537 5960 9571
rect 5908 9528 5960 9537
rect 6368 9528 6420 9580
rect 11980 9571 12032 9580
rect 11980 9537 11989 9571
rect 11989 9537 12023 9571
rect 12023 9537 12032 9571
rect 11980 9528 12032 9537
rect 14188 9460 14240 9512
rect 16672 9503 16724 9512
rect 16672 9469 16681 9503
rect 16681 9469 16715 9503
rect 16715 9469 16724 9503
rect 16672 9460 16724 9469
rect 16948 9503 17000 9512
rect 16948 9469 16957 9503
rect 16957 9469 16991 9503
rect 16991 9469 17000 9503
rect 16948 9460 17000 9469
rect 2688 9324 2740 9376
rect 4252 9324 4304 9376
rect 5632 9367 5684 9376
rect 5632 9333 5641 9367
rect 5641 9333 5675 9367
rect 5675 9333 5684 9367
rect 5632 9324 5684 9333
rect 14188 9324 14240 9376
rect 17960 9324 18012 9376
rect 18328 9324 18380 9376
rect 2350 9222 2402 9274
rect 2414 9222 2466 9274
rect 2478 9222 2530 9274
rect 2542 9222 2594 9274
rect 2606 9222 2658 9274
rect 2872 9120 2924 9172
rect 17408 9120 17460 9172
rect 18788 9163 18840 9172
rect 18788 9129 18797 9163
rect 18797 9129 18831 9163
rect 18831 9129 18840 9163
rect 18788 9120 18840 9129
rect 848 9052 900 9104
rect 1860 8916 1912 8968
rect 5632 8984 5684 9036
rect 8300 8984 8352 9036
rect 2136 8916 2188 8968
rect 5816 8916 5868 8968
rect 8576 8916 8628 8968
rect 9128 8959 9180 8968
rect 9128 8925 9137 8959
rect 9137 8925 9171 8959
rect 9171 8925 9180 8959
rect 9128 8916 9180 8925
rect 9312 8959 9364 8968
rect 9312 8925 9321 8959
rect 9321 8925 9355 8959
rect 9355 8925 9364 8959
rect 9312 8916 9364 8925
rect 13728 8916 13780 8968
rect 14188 8959 14240 8968
rect 14188 8925 14197 8959
rect 14197 8925 14231 8959
rect 14231 8925 14240 8959
rect 14188 8916 14240 8925
rect 16580 8916 16632 8968
rect 18328 8959 18380 8968
rect 18328 8925 18337 8959
rect 18337 8925 18371 8959
rect 18371 8925 18380 8959
rect 18328 8916 18380 8925
rect 18604 8959 18656 8968
rect 18604 8925 18613 8959
rect 18613 8925 18647 8959
rect 18647 8925 18656 8959
rect 18604 8916 18656 8925
rect 9864 8848 9916 8900
rect 9680 8780 9732 8832
rect 9772 8780 9824 8832
rect 11980 8780 12032 8832
rect 15384 8780 15436 8832
rect 16028 8780 16080 8832
rect 18512 8823 18564 8832
rect 18512 8789 18521 8823
rect 18521 8789 18555 8823
rect 18555 8789 18564 8823
rect 18512 8780 18564 8789
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 2688 8576 2740 8628
rect 9128 8576 9180 8628
rect 2228 8508 2280 8560
rect 5816 8508 5868 8560
rect 17408 8508 17460 8560
rect 4252 8483 4304 8492
rect 4252 8449 4261 8483
rect 4261 8449 4295 8483
rect 4295 8449 4304 8483
rect 4252 8440 4304 8449
rect 4620 8483 4672 8492
rect 4620 8449 4629 8483
rect 4629 8449 4663 8483
rect 4663 8449 4672 8483
rect 4620 8440 4672 8449
rect 8116 8483 8168 8492
rect 8116 8449 8125 8483
rect 8125 8449 8159 8483
rect 8159 8449 8168 8483
rect 8116 8440 8168 8449
rect 9312 8440 9364 8492
rect 9772 8483 9824 8492
rect 9772 8449 9781 8483
rect 9781 8449 9815 8483
rect 9815 8449 9824 8483
rect 9772 8440 9824 8449
rect 9864 8440 9916 8492
rect 14188 8440 14240 8492
rect 16672 8440 16724 8492
rect 18236 8440 18288 8492
rect 2872 8415 2924 8424
rect 2872 8381 2881 8415
rect 2881 8381 2915 8415
rect 2915 8381 2924 8415
rect 2872 8372 2924 8381
rect 15660 8372 15712 8424
rect 15752 8415 15804 8424
rect 15752 8381 15761 8415
rect 15761 8381 15795 8415
rect 15795 8381 15804 8415
rect 15752 8372 15804 8381
rect 17132 8415 17184 8424
rect 17132 8381 17141 8415
rect 17141 8381 17175 8415
rect 17175 8381 17184 8415
rect 17132 8372 17184 8381
rect 4160 8304 4212 8356
rect 4252 8304 4304 8356
rect 1768 8236 1820 8288
rect 18144 8236 18196 8288
rect 2350 8134 2402 8186
rect 2414 8134 2466 8186
rect 2478 8134 2530 8186
rect 2542 8134 2594 8186
rect 2606 8134 2658 8186
rect 1308 8032 1360 8084
rect 2228 8032 2280 8084
rect 1768 7828 1820 7880
rect 1860 7803 1912 7812
rect 1860 7769 1869 7803
rect 1869 7769 1903 7803
rect 1903 7769 1912 7803
rect 1860 7760 1912 7769
rect 2136 7828 2188 7880
rect 2596 7828 2648 7880
rect 3608 7828 3660 7880
rect 8576 8032 8628 8084
rect 15752 8032 15804 8084
rect 17132 8032 17184 8084
rect 18236 8032 18288 8084
rect 4160 8007 4212 8016
rect 4160 7973 4169 8007
rect 4169 7973 4203 8007
rect 4203 7973 4212 8007
rect 4160 7964 4212 7973
rect 3884 7939 3936 7948
rect 3884 7905 3893 7939
rect 3893 7905 3927 7939
rect 3927 7905 3936 7939
rect 3884 7896 3936 7905
rect 3976 7939 4028 7948
rect 3976 7905 3985 7939
rect 3985 7905 4019 7939
rect 4019 7905 4028 7939
rect 3976 7896 4028 7905
rect 5816 7896 5868 7948
rect 14096 7939 14148 7948
rect 14096 7905 14105 7939
rect 14105 7905 14139 7939
rect 14139 7905 14148 7939
rect 14096 7896 14148 7905
rect 15384 7896 15436 7948
rect 6828 7828 6880 7880
rect 9128 7871 9180 7880
rect 9128 7837 9137 7871
rect 9137 7837 9171 7871
rect 9171 7837 9180 7871
rect 9128 7828 9180 7837
rect 13452 7828 13504 7880
rect 13728 7871 13780 7880
rect 13728 7837 13737 7871
rect 13737 7837 13771 7871
rect 13771 7837 13780 7871
rect 13728 7828 13780 7837
rect 15936 7871 15988 7880
rect 15936 7837 15945 7871
rect 15945 7837 15979 7871
rect 15979 7837 15988 7871
rect 15936 7828 15988 7837
rect 16028 7871 16080 7880
rect 16028 7837 16038 7871
rect 16038 7837 16072 7871
rect 16072 7837 16080 7871
rect 16028 7828 16080 7837
rect 17408 7871 17460 7880
rect 17408 7837 17417 7871
rect 17417 7837 17451 7871
rect 17451 7837 17460 7871
rect 17408 7828 17460 7837
rect 5540 7760 5592 7812
rect 14648 7760 14700 7812
rect 17684 7871 17736 7880
rect 17684 7837 17693 7871
rect 17693 7837 17727 7871
rect 17727 7837 17736 7871
rect 17684 7828 17736 7837
rect 18052 7871 18104 7880
rect 18052 7837 18060 7871
rect 18060 7837 18094 7871
rect 18094 7837 18104 7871
rect 18052 7828 18104 7837
rect 18144 7871 18196 7880
rect 18144 7837 18153 7871
rect 18153 7837 18187 7871
rect 18187 7837 18196 7871
rect 18144 7828 18196 7837
rect 2504 7735 2556 7744
rect 2504 7701 2513 7735
rect 2513 7701 2547 7735
rect 2547 7701 2556 7735
rect 2504 7692 2556 7701
rect 4804 7692 4856 7744
rect 9036 7735 9088 7744
rect 9036 7701 9045 7735
rect 9045 7701 9079 7735
rect 9079 7701 9088 7735
rect 9036 7692 9088 7701
rect 15752 7692 15804 7744
rect 16580 7692 16632 7744
rect 18604 7871 18656 7880
rect 18604 7837 18613 7871
rect 18613 7837 18647 7871
rect 18647 7837 18656 7871
rect 18604 7828 18656 7837
rect 18788 7735 18840 7744
rect 18788 7701 18797 7735
rect 18797 7701 18831 7735
rect 18831 7701 18840 7735
rect 18788 7692 18840 7701
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 1308 7488 1360 7540
rect 2872 7488 2924 7540
rect 3884 7488 3936 7540
rect 5540 7488 5592 7540
rect 5908 7488 5960 7540
rect 6828 7488 6880 7540
rect 4620 7420 4672 7472
rect 2504 7352 2556 7404
rect 3700 7395 3752 7404
rect 3700 7361 3709 7395
rect 3709 7361 3743 7395
rect 3743 7361 3752 7395
rect 3700 7352 3752 7361
rect 3884 7352 3936 7404
rect 4252 7395 4304 7404
rect 4252 7361 4261 7395
rect 4261 7361 4295 7395
rect 4295 7361 4304 7395
rect 4252 7352 4304 7361
rect 4528 7395 4580 7404
rect 4528 7361 4537 7395
rect 4537 7361 4571 7395
rect 4571 7361 4580 7395
rect 4528 7352 4580 7361
rect 4804 7395 4856 7404
rect 4804 7361 4813 7395
rect 4813 7361 4847 7395
rect 4847 7361 4856 7395
rect 4804 7352 4856 7361
rect 5908 7352 5960 7404
rect 3792 7216 3844 7268
rect 4252 7216 4304 7268
rect 6000 7216 6052 7268
rect 7288 7352 7340 7404
rect 14648 7531 14700 7540
rect 14648 7497 14657 7531
rect 14657 7497 14691 7531
rect 14691 7497 14700 7531
rect 14648 7488 14700 7497
rect 15292 7488 15344 7540
rect 17684 7488 17736 7540
rect 8300 7420 8352 7472
rect 9036 7420 9088 7472
rect 13728 7352 13780 7404
rect 15752 7420 15804 7472
rect 17408 7420 17460 7472
rect 7564 7284 7616 7336
rect 9588 7327 9640 7336
rect 9588 7293 9597 7327
rect 9597 7293 9631 7327
rect 9631 7293 9640 7327
rect 9588 7284 9640 7293
rect 9772 7327 9824 7336
rect 9772 7293 9781 7327
rect 9781 7293 9815 7327
rect 9815 7293 9824 7327
rect 9772 7284 9824 7293
rect 15292 7352 15344 7404
rect 15384 7395 15436 7404
rect 15384 7361 15393 7395
rect 15393 7361 15427 7395
rect 15427 7361 15436 7395
rect 15384 7352 15436 7361
rect 15476 7395 15528 7404
rect 15476 7361 15485 7395
rect 15485 7361 15519 7395
rect 15519 7361 15528 7395
rect 15476 7352 15528 7361
rect 16028 7352 16080 7404
rect 18144 7395 18196 7404
rect 18144 7361 18153 7395
rect 18153 7361 18187 7395
rect 18187 7361 18196 7395
rect 18144 7352 18196 7361
rect 18328 7352 18380 7404
rect 15844 7284 15896 7336
rect 6828 7216 6880 7268
rect 4068 7191 4120 7200
rect 4068 7157 4077 7191
rect 4077 7157 4111 7191
rect 4111 7157 4120 7191
rect 4068 7148 4120 7157
rect 6368 7191 6420 7200
rect 6368 7157 6377 7191
rect 6377 7157 6411 7191
rect 6411 7157 6420 7191
rect 6368 7148 6420 7157
rect 7104 7148 7156 7200
rect 9496 7191 9548 7200
rect 9496 7157 9505 7191
rect 9505 7157 9539 7191
rect 9539 7157 9548 7191
rect 9496 7148 9548 7157
rect 9680 7148 9732 7200
rect 15384 7148 15436 7200
rect 18512 7148 18564 7200
rect 18788 7191 18840 7200
rect 18788 7157 18797 7191
rect 18797 7157 18831 7191
rect 18831 7157 18840 7191
rect 18788 7148 18840 7157
rect 2350 7046 2402 7098
rect 2414 7046 2466 7098
rect 2478 7046 2530 7098
rect 2542 7046 2594 7098
rect 2606 7046 2658 7098
rect 3976 6987 4028 6996
rect 3976 6953 3985 6987
rect 3985 6953 4019 6987
rect 4019 6953 4028 6987
rect 3976 6944 4028 6953
rect 6368 6944 6420 6996
rect 7288 6987 7340 6996
rect 7288 6953 7297 6987
rect 7297 6953 7331 6987
rect 7331 6953 7340 6987
rect 7288 6944 7340 6953
rect 15844 6987 15896 6996
rect 15844 6953 15874 6987
rect 15874 6953 15896 6987
rect 15844 6944 15896 6953
rect 18328 6987 18380 6996
rect 18328 6953 18337 6987
rect 18337 6953 18371 6987
rect 18371 6953 18380 6987
rect 18328 6944 18380 6953
rect 18604 6987 18656 6996
rect 18604 6953 18613 6987
rect 18613 6953 18647 6987
rect 18647 6953 18656 6987
rect 18604 6944 18656 6953
rect 9772 6876 9824 6928
rect 3700 6808 3752 6860
rect 4068 6851 4120 6860
rect 4068 6817 4077 6851
rect 4077 6817 4111 6851
rect 4111 6817 4120 6851
rect 4068 6808 4120 6817
rect 5816 6808 5868 6860
rect 14096 6808 14148 6860
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 3792 6783 3844 6792
rect 3792 6749 3801 6783
rect 3801 6749 3835 6783
rect 3835 6749 3844 6783
rect 3792 6740 3844 6749
rect 3884 6783 3936 6792
rect 3884 6749 3893 6783
rect 3893 6749 3927 6783
rect 3927 6749 3936 6783
rect 3884 6740 3936 6749
rect 3976 6740 4028 6792
rect 8300 6740 8352 6792
rect 8576 6783 8628 6792
rect 8576 6749 8585 6783
rect 8585 6749 8619 6783
rect 8619 6749 8628 6783
rect 8576 6740 8628 6749
rect 9036 6783 9088 6792
rect 9036 6749 9045 6783
rect 9045 6749 9079 6783
rect 9079 6749 9088 6783
rect 9036 6740 9088 6749
rect 9496 6740 9548 6792
rect 14372 6740 14424 6792
rect 14648 6740 14700 6792
rect 16580 6808 16632 6860
rect 17224 6808 17276 6860
rect 15568 6783 15620 6792
rect 15568 6749 15577 6783
rect 15577 6749 15611 6783
rect 15611 6749 15620 6783
rect 15568 6740 15620 6749
rect 18604 6740 18656 6792
rect 1676 6715 1728 6724
rect 1676 6681 1685 6715
rect 1685 6681 1719 6715
rect 1719 6681 1728 6715
rect 1676 6672 1728 6681
rect 2412 6672 2464 6724
rect 7104 6672 7156 6724
rect 3424 6604 3476 6656
rect 9312 6604 9364 6656
rect 16856 6672 16908 6724
rect 14464 6647 14516 6656
rect 14464 6613 14473 6647
rect 14473 6613 14507 6647
rect 14507 6613 14516 6647
rect 14464 6604 14516 6613
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 2412 6443 2464 6452
rect 2412 6409 2421 6443
rect 2421 6409 2455 6443
rect 2455 6409 2464 6443
rect 2412 6400 2464 6409
rect 3976 6400 4028 6452
rect 9588 6400 9640 6452
rect 14464 6443 14516 6452
rect 14464 6409 14473 6443
rect 14473 6409 14507 6443
rect 14507 6409 14516 6443
rect 14464 6400 14516 6409
rect 14556 6400 14608 6452
rect 16856 6400 16908 6452
rect 18052 6400 18104 6452
rect 12532 6375 12584 6384
rect 12532 6341 12541 6375
rect 12541 6341 12575 6375
rect 12575 6341 12584 6375
rect 12532 6332 12584 6341
rect 848 6264 900 6316
rect 1584 6264 1636 6316
rect 2136 6264 2188 6316
rect 2688 6264 2740 6316
rect 2780 6264 2832 6316
rect 3700 6264 3752 6316
rect 9128 6264 9180 6316
rect 9772 6264 9824 6316
rect 15292 6332 15344 6384
rect 16580 6332 16632 6384
rect 16948 6332 17000 6384
rect 14556 6307 14608 6316
rect 14556 6273 14565 6307
rect 14565 6273 14599 6307
rect 14599 6273 14608 6307
rect 14556 6264 14608 6273
rect 14648 6264 14700 6316
rect 17224 6264 17276 6316
rect 17868 6264 17920 6316
rect 18604 6264 18656 6316
rect 18788 6307 18840 6316
rect 18788 6273 18797 6307
rect 18797 6273 18831 6307
rect 18831 6273 18840 6307
rect 18788 6264 18840 6273
rect 1676 6171 1728 6180
rect 1676 6137 1685 6171
rect 1685 6137 1719 6171
rect 1719 6137 1728 6171
rect 1676 6128 1728 6137
rect 2228 6128 2280 6180
rect 3424 6196 3476 6248
rect 6920 6196 6972 6248
rect 7564 6239 7616 6248
rect 7564 6205 7573 6239
rect 7573 6205 7607 6239
rect 7607 6205 7616 6239
rect 7564 6196 7616 6205
rect 8852 6196 8904 6248
rect 15016 6239 15068 6248
rect 15016 6205 15025 6239
rect 15025 6205 15059 6239
rect 15059 6205 15068 6239
rect 15016 6196 15068 6205
rect 17500 6128 17552 6180
rect 1952 6103 2004 6112
rect 1952 6069 1961 6103
rect 1961 6069 1995 6103
rect 1995 6069 2004 6103
rect 1952 6060 2004 6069
rect 13728 6060 13780 6112
rect 17316 6060 17368 6112
rect 2350 5958 2402 6010
rect 2414 5958 2466 6010
rect 2478 5958 2530 6010
rect 2542 5958 2594 6010
rect 2606 5958 2658 6010
rect 2320 5856 2372 5908
rect 3976 5856 4028 5908
rect 8300 5856 8352 5908
rect 8852 5856 8904 5908
rect 14556 5856 14608 5908
rect 2780 5788 2832 5840
rect 3700 5788 3752 5840
rect 1400 5720 1452 5772
rect 2688 5720 2740 5772
rect 8024 5788 8076 5840
rect 6828 5720 6880 5772
rect 1492 5516 1544 5568
rect 1768 5516 1820 5568
rect 2228 5652 2280 5704
rect 2320 5695 2372 5704
rect 2320 5661 2329 5695
rect 2329 5661 2363 5695
rect 2363 5661 2372 5695
rect 2320 5652 2372 5661
rect 3516 5652 3568 5704
rect 3792 5695 3844 5704
rect 3792 5661 3801 5695
rect 3801 5661 3835 5695
rect 3835 5661 3844 5695
rect 3792 5652 3844 5661
rect 3976 5695 4028 5704
rect 3976 5661 3985 5695
rect 3985 5661 4019 5695
rect 4019 5661 4028 5695
rect 3976 5652 4028 5661
rect 5908 5652 5960 5704
rect 7012 5652 7064 5704
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 8760 5695 8812 5704
rect 8760 5661 8769 5695
rect 8769 5661 8803 5695
rect 8803 5661 8812 5695
rect 8760 5652 8812 5661
rect 10968 5788 11020 5840
rect 9220 5720 9272 5772
rect 11888 5720 11940 5772
rect 9312 5695 9364 5704
rect 9312 5661 9321 5695
rect 9321 5661 9355 5695
rect 9355 5661 9364 5695
rect 9312 5652 9364 5661
rect 9588 5652 9640 5704
rect 9772 5652 9824 5704
rect 10968 5652 11020 5704
rect 13728 5788 13780 5840
rect 16028 5831 16080 5840
rect 16028 5797 16037 5831
rect 16037 5797 16071 5831
rect 16071 5797 16080 5831
rect 16028 5788 16080 5797
rect 16580 5899 16632 5908
rect 16580 5865 16589 5899
rect 16589 5865 16623 5899
rect 16623 5865 16632 5899
rect 16580 5856 16632 5865
rect 18604 5899 18656 5908
rect 18604 5865 18613 5899
rect 18613 5865 18647 5899
rect 18647 5865 18656 5899
rect 18604 5856 18656 5865
rect 15568 5720 15620 5772
rect 17868 5720 17920 5772
rect 3608 5584 3660 5636
rect 13452 5652 13504 5704
rect 14280 5652 14332 5704
rect 13268 5584 13320 5636
rect 17132 5627 17184 5636
rect 17132 5593 17141 5627
rect 17141 5593 17175 5627
rect 17175 5593 17184 5627
rect 17132 5584 17184 5593
rect 18144 5584 18196 5636
rect 2780 5516 2832 5568
rect 5816 5559 5868 5568
rect 5816 5525 5825 5559
rect 5825 5525 5859 5559
rect 5859 5525 5868 5559
rect 5816 5516 5868 5525
rect 6920 5516 6972 5568
rect 8576 5516 8628 5568
rect 10968 5559 11020 5568
rect 10968 5525 10977 5559
rect 10977 5525 11011 5559
rect 11011 5525 11020 5559
rect 10968 5516 11020 5525
rect 12072 5559 12124 5568
rect 12072 5525 12081 5559
rect 12081 5525 12115 5559
rect 12115 5525 12124 5559
rect 12072 5516 12124 5525
rect 12532 5516 12584 5568
rect 14740 5516 14792 5568
rect 16488 5516 16540 5568
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 2780 5312 2832 5364
rect 3516 5355 3568 5364
rect 3516 5321 3525 5355
rect 3525 5321 3559 5355
rect 3559 5321 3568 5355
rect 3516 5312 3568 5321
rect 1768 5287 1820 5296
rect 1768 5253 1777 5287
rect 1777 5253 1811 5287
rect 1811 5253 1820 5287
rect 1768 5244 1820 5253
rect 3976 5244 4028 5296
rect 1400 5176 1452 5228
rect 2872 5176 2924 5228
rect 3608 5219 3660 5228
rect 3608 5185 3617 5219
rect 3617 5185 3651 5219
rect 3651 5185 3660 5219
rect 3608 5176 3660 5185
rect 3792 5219 3844 5228
rect 3792 5185 3801 5219
rect 3801 5185 3835 5219
rect 3835 5185 3844 5219
rect 3792 5176 3844 5185
rect 5816 5312 5868 5364
rect 6000 5287 6052 5296
rect 6000 5253 6009 5287
rect 6009 5253 6043 5287
rect 6043 5253 6052 5287
rect 6000 5244 6052 5253
rect 9036 5312 9088 5364
rect 11244 5312 11296 5364
rect 13268 5355 13320 5364
rect 13268 5321 13277 5355
rect 13277 5321 13311 5355
rect 13311 5321 13320 5355
rect 13268 5312 13320 5321
rect 15016 5355 15068 5364
rect 15016 5321 15025 5355
rect 15025 5321 15059 5355
rect 15059 5321 15068 5355
rect 15016 5312 15068 5321
rect 17132 5312 17184 5364
rect 18144 5312 18196 5364
rect 18788 5355 18840 5364
rect 18788 5321 18797 5355
rect 18797 5321 18831 5355
rect 18831 5321 18840 5355
rect 18788 5312 18840 5321
rect 2228 5108 2280 5160
rect 4068 5040 4120 5092
rect 5356 5151 5408 5160
rect 5356 5117 5365 5151
rect 5365 5117 5399 5151
rect 5399 5117 5408 5151
rect 5356 5108 5408 5117
rect 7012 5219 7064 5228
rect 7012 5185 7021 5219
rect 7021 5185 7055 5219
rect 7055 5185 7064 5219
rect 7012 5176 7064 5185
rect 8024 5287 8076 5296
rect 8024 5253 8033 5287
rect 8033 5253 8067 5287
rect 8067 5253 8076 5287
rect 8024 5244 8076 5253
rect 9588 5244 9640 5296
rect 10968 5244 11020 5296
rect 11428 5244 11480 5296
rect 12532 5244 12584 5296
rect 14280 5244 14332 5296
rect 7656 5176 7708 5228
rect 6920 5108 6972 5160
rect 11060 5151 11112 5160
rect 11060 5117 11069 5151
rect 11069 5117 11103 5151
rect 11103 5117 11112 5151
rect 11060 5108 11112 5117
rect 11520 5151 11572 5160
rect 11520 5117 11529 5151
rect 11529 5117 11563 5151
rect 11563 5117 11572 5151
rect 11520 5108 11572 5117
rect 14740 5219 14792 5228
rect 14740 5185 14750 5219
rect 14750 5185 14784 5219
rect 14784 5185 14792 5219
rect 17224 5244 17276 5296
rect 14740 5176 14792 5185
rect 15936 5108 15988 5160
rect 17132 5176 17184 5228
rect 17224 5108 17276 5160
rect 17316 5040 17368 5092
rect 17500 5219 17552 5228
rect 17500 5185 17509 5219
rect 17509 5185 17543 5219
rect 17543 5185 17552 5219
rect 17500 5176 17552 5185
rect 17684 5219 17736 5228
rect 17684 5185 17693 5219
rect 17693 5185 17727 5219
rect 17727 5185 17736 5219
rect 17684 5176 17736 5185
rect 18512 5176 18564 5228
rect 18144 5040 18196 5092
rect 7012 4972 7064 5024
rect 7472 5015 7524 5024
rect 7472 4981 7481 5015
rect 7481 4981 7515 5015
rect 7515 4981 7524 5015
rect 7472 4972 7524 4981
rect 10692 4972 10744 5024
rect 15384 4972 15436 5024
rect 17132 4972 17184 5024
rect 17868 4972 17920 5024
rect 18052 4972 18104 5024
rect 2350 4870 2402 4922
rect 2414 4870 2466 4922
rect 2478 4870 2530 4922
rect 2542 4870 2594 4922
rect 2606 4870 2658 4922
rect 2872 4768 2924 4820
rect 3792 4768 3844 4820
rect 7656 4768 7708 4820
rect 9588 4811 9640 4820
rect 9588 4777 9597 4811
rect 9597 4777 9631 4811
rect 9631 4777 9640 4811
rect 9588 4768 9640 4777
rect 11060 4768 11112 4820
rect 16396 4811 16448 4820
rect 16396 4777 16405 4811
rect 16405 4777 16439 4811
rect 16439 4777 16448 4811
rect 16396 4768 16448 4777
rect 1952 4632 2004 4684
rect 848 4564 900 4616
rect 2136 4564 2188 4616
rect 3608 4632 3660 4684
rect 3700 4564 3752 4616
rect 5356 4564 5408 4616
rect 5540 4564 5592 4616
rect 6920 4632 6972 4684
rect 12072 4632 12124 4684
rect 9772 4564 9824 4616
rect 10692 4607 10744 4616
rect 10692 4573 10701 4607
rect 10701 4573 10735 4607
rect 10735 4573 10744 4607
rect 10692 4564 10744 4573
rect 11152 4564 11204 4616
rect 2044 4496 2096 4548
rect 4160 4471 4212 4480
rect 4160 4437 4169 4471
rect 4169 4437 4203 4471
rect 4203 4437 4212 4471
rect 4160 4428 4212 4437
rect 7012 4496 7064 4548
rect 8668 4496 8720 4548
rect 11428 4607 11480 4616
rect 11428 4573 11437 4607
rect 11437 4573 11471 4607
rect 11471 4573 11480 4607
rect 11428 4564 11480 4573
rect 13728 4564 13780 4616
rect 15936 4564 15988 4616
rect 17776 4564 17828 4616
rect 18236 4607 18288 4616
rect 18236 4573 18245 4607
rect 18245 4573 18279 4607
rect 18279 4573 18288 4607
rect 18236 4564 18288 4573
rect 18328 4564 18380 4616
rect 11336 4496 11388 4548
rect 6644 4428 6696 4480
rect 12624 4471 12676 4480
rect 12624 4437 12633 4471
rect 12633 4437 12667 4471
rect 12667 4437 12676 4471
rect 12624 4428 12676 4437
rect 15384 4496 15436 4548
rect 16580 4428 16632 4480
rect 17684 4428 17736 4480
rect 18788 4471 18840 4480
rect 18788 4437 18797 4471
rect 18797 4437 18831 4471
rect 18831 4437 18840 4471
rect 18788 4428 18840 4437
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 4160 4224 4212 4276
rect 5356 4224 5408 4276
rect 11336 4224 11388 4276
rect 1676 4131 1728 4140
rect 1676 4097 1685 4131
rect 1685 4097 1719 4131
rect 1719 4097 1728 4131
rect 1676 4088 1728 4097
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 1952 4020 2004 4072
rect 2228 4156 2280 4208
rect 3240 4131 3292 4140
rect 3240 4097 3249 4131
rect 3249 4097 3283 4131
rect 3283 4097 3292 4131
rect 3240 4088 3292 4097
rect 5724 4088 5776 4140
rect 8116 4156 8168 4208
rect 6644 4131 6696 4140
rect 6644 4097 6653 4131
rect 6653 4097 6687 4131
rect 6687 4097 6696 4131
rect 6644 4088 6696 4097
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 2688 4020 2740 4072
rect 7104 4088 7156 4140
rect 7472 4088 7524 4140
rect 8852 4131 8904 4140
rect 8852 4097 8891 4131
rect 8891 4097 8904 4131
rect 8852 4088 8904 4097
rect 10692 4088 10744 4140
rect 11888 4088 11940 4140
rect 7288 4020 7340 4072
rect 11980 4020 12032 4072
rect 12624 4131 12676 4140
rect 12624 4097 12633 4131
rect 12633 4097 12667 4131
rect 12667 4097 12676 4131
rect 12624 4088 12676 4097
rect 12992 4088 13044 4140
rect 13452 4131 13504 4140
rect 13452 4097 13461 4131
rect 13461 4097 13495 4131
rect 13495 4097 13504 4131
rect 13452 4088 13504 4097
rect 15200 4131 15252 4140
rect 15200 4097 15209 4131
rect 15209 4097 15243 4131
rect 15243 4097 15252 4131
rect 15200 4088 15252 4097
rect 8300 3952 8352 4004
rect 12900 3952 12952 4004
rect 16396 4088 16448 4140
rect 18420 4088 18472 4140
rect 15844 4063 15896 4072
rect 15844 4029 15853 4063
rect 15853 4029 15887 4063
rect 15887 4029 15896 4063
rect 15844 4020 15896 4029
rect 17040 4063 17092 4072
rect 17040 4029 17049 4063
rect 17049 4029 17083 4063
rect 17083 4029 17092 4063
rect 17040 4020 17092 4029
rect 17316 4063 17368 4072
rect 17316 4029 17325 4063
rect 17325 4029 17359 4063
rect 17359 4029 17368 4063
rect 17316 4020 17368 4029
rect 15936 3952 15988 4004
rect 5816 3884 5868 3936
rect 7104 3927 7156 3936
rect 7104 3893 7113 3927
rect 7113 3893 7147 3927
rect 7147 3893 7156 3927
rect 7104 3884 7156 3893
rect 8392 3884 8444 3936
rect 12256 3927 12308 3936
rect 12256 3893 12265 3927
rect 12265 3893 12299 3927
rect 12299 3893 12308 3927
rect 12256 3884 12308 3893
rect 13452 3884 13504 3936
rect 14372 3884 14424 3936
rect 17500 3884 17552 3936
rect 18788 3927 18840 3936
rect 18788 3893 18797 3927
rect 18797 3893 18831 3927
rect 18831 3893 18840 3927
rect 18788 3884 18840 3893
rect 2350 3782 2402 3834
rect 2414 3782 2466 3834
rect 2478 3782 2530 3834
rect 2542 3782 2594 3834
rect 2606 3782 2658 3834
rect 2136 3680 2188 3732
rect 6828 3680 6880 3732
rect 10692 3723 10744 3732
rect 10692 3689 10701 3723
rect 10701 3689 10735 3723
rect 10735 3689 10744 3723
rect 10692 3680 10744 3689
rect 11888 3723 11940 3732
rect 11888 3689 11897 3723
rect 11897 3689 11931 3723
rect 11931 3689 11940 3723
rect 11888 3680 11940 3689
rect 12256 3680 12308 3732
rect 12992 3680 13044 3732
rect 6920 3612 6972 3664
rect 15844 3723 15896 3732
rect 15844 3689 15853 3723
rect 15853 3689 15887 3723
rect 15887 3689 15896 3723
rect 15844 3680 15896 3689
rect 15936 3680 15988 3732
rect 17316 3680 17368 3732
rect 18328 3723 18380 3732
rect 18328 3689 18337 3723
rect 18337 3689 18371 3723
rect 18371 3689 18380 3723
rect 18328 3680 18380 3689
rect 18420 3680 18472 3732
rect 2688 3544 2740 3596
rect 5540 3587 5592 3596
rect 5540 3553 5549 3587
rect 5549 3553 5583 3587
rect 5583 3553 5592 3587
rect 5540 3544 5592 3553
rect 5816 3587 5868 3596
rect 5816 3553 5825 3587
rect 5825 3553 5859 3587
rect 5859 3553 5868 3587
rect 5816 3544 5868 3553
rect 7288 3587 7340 3596
rect 7288 3553 7297 3587
rect 7297 3553 7331 3587
rect 7331 3553 7340 3587
rect 7288 3544 7340 3553
rect 848 3476 900 3528
rect 3240 3476 3292 3528
rect 8668 3544 8720 3596
rect 11520 3544 11572 3596
rect 13728 3544 13780 3596
rect 7104 3408 7156 3460
rect 8300 3519 8352 3528
rect 8300 3485 8309 3519
rect 8309 3485 8343 3519
rect 8343 3485 8352 3519
rect 8300 3476 8352 3485
rect 8392 3519 8444 3528
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 8392 3476 8444 3485
rect 8852 3476 8904 3528
rect 11428 3476 11480 3528
rect 11888 3519 11940 3528
rect 11888 3485 11927 3519
rect 11927 3485 11940 3519
rect 11888 3476 11940 3485
rect 3976 3340 4028 3392
rect 6828 3340 6880 3392
rect 9772 3408 9824 3460
rect 13452 3408 13504 3460
rect 13728 3340 13780 3392
rect 17868 3612 17920 3664
rect 16580 3476 16632 3528
rect 17776 3544 17828 3596
rect 17592 3519 17644 3528
rect 17592 3485 17601 3519
rect 17601 3485 17635 3519
rect 17635 3485 17644 3519
rect 17592 3476 17644 3485
rect 17684 3519 17736 3528
rect 17684 3485 17693 3519
rect 17693 3485 17727 3519
rect 17727 3485 17736 3519
rect 17684 3476 17736 3485
rect 17868 3519 17920 3528
rect 17868 3485 17877 3519
rect 17877 3485 17911 3519
rect 17911 3485 17920 3519
rect 17868 3476 17920 3485
rect 18236 3544 18288 3596
rect 18788 3544 18840 3596
rect 14372 3451 14424 3460
rect 14372 3417 14381 3451
rect 14381 3417 14415 3451
rect 14415 3417 14424 3451
rect 14372 3408 14424 3417
rect 15844 3408 15896 3460
rect 16672 3408 16724 3460
rect 17224 3408 17276 3460
rect 17040 3340 17092 3392
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 1676 3136 1728 3188
rect 3976 3111 4028 3120
rect 3976 3077 3985 3111
rect 3985 3077 4019 3111
rect 4019 3077 4028 3111
rect 3976 3068 4028 3077
rect 848 3000 900 3052
rect 2688 3000 2740 3052
rect 5724 3043 5776 3052
rect 5724 3009 5733 3043
rect 5733 3009 5767 3043
rect 5767 3009 5776 3043
rect 5724 3000 5776 3009
rect 8760 3136 8812 3188
rect 7012 3068 7064 3120
rect 8392 3068 8444 3120
rect 6920 3000 6972 3052
rect 6644 2864 6696 2916
rect 9772 3179 9824 3188
rect 9772 3145 9781 3179
rect 9781 3145 9815 3179
rect 9815 3145 9824 3179
rect 9772 3136 9824 3145
rect 9864 3136 9916 3188
rect 11704 3136 11756 3188
rect 15200 3136 15252 3188
rect 10968 3068 11020 3120
rect 9864 3000 9916 3052
rect 10692 3000 10744 3052
rect 12072 3068 12124 3120
rect 12532 3068 12584 3120
rect 15476 3111 15528 3120
rect 15476 3077 15485 3111
rect 15485 3077 15519 3111
rect 15519 3077 15528 3111
rect 15476 3068 15528 3077
rect 15844 3179 15896 3188
rect 15844 3145 15853 3179
rect 15853 3145 15887 3179
rect 15887 3145 15896 3179
rect 15844 3136 15896 3145
rect 16948 3136 17000 3188
rect 11244 3000 11296 3052
rect 11520 3043 11572 3052
rect 11520 3009 11529 3043
rect 11529 3009 11563 3043
rect 11563 3009 11572 3043
rect 11520 3000 11572 3009
rect 11888 2932 11940 2984
rect 12440 2932 12492 2984
rect 13728 3043 13780 3052
rect 13728 3009 13737 3043
rect 13737 3009 13771 3043
rect 13771 3009 13780 3043
rect 13728 3000 13780 3009
rect 17040 3068 17092 3120
rect 17224 3068 17276 3120
rect 11152 2864 11204 2916
rect 6736 2796 6788 2848
rect 6828 2839 6880 2848
rect 6828 2805 6837 2839
rect 6837 2805 6871 2839
rect 6871 2805 6880 2839
rect 6828 2796 6880 2805
rect 9312 2796 9364 2848
rect 10600 2796 10652 2848
rect 11428 2864 11480 2916
rect 16028 2932 16080 2984
rect 16948 2975 17000 2984
rect 16948 2941 16957 2975
rect 16957 2941 16991 2975
rect 16991 2941 17000 2975
rect 16948 2932 17000 2941
rect 12164 2796 12216 2848
rect 12256 2796 12308 2848
rect 13820 2796 13872 2848
rect 14464 2796 14516 2848
rect 16672 2864 16724 2916
rect 16580 2796 16632 2848
rect 18604 2796 18656 2848
rect 2350 2694 2402 2746
rect 2414 2694 2466 2746
rect 2478 2694 2530 2746
rect 2542 2694 2594 2746
rect 2606 2694 2658 2746
rect 6828 2592 6880 2644
rect 7012 2592 7064 2644
rect 8392 2592 8444 2644
rect 11060 2635 11112 2644
rect 11060 2601 11069 2635
rect 11069 2601 11103 2635
rect 11103 2601 11112 2635
rect 11060 2592 11112 2601
rect 12532 2592 12584 2644
rect 15476 2592 15528 2644
rect 17224 2592 17276 2644
rect 17408 2592 17460 2644
rect 17776 2635 17828 2644
rect 17776 2601 17785 2635
rect 17785 2601 17819 2635
rect 17819 2601 17828 2635
rect 17776 2592 17828 2601
rect 18052 2635 18104 2644
rect 18052 2601 18061 2635
rect 18061 2601 18095 2635
rect 18095 2601 18104 2635
rect 18052 2592 18104 2601
rect 18788 2635 18840 2644
rect 18788 2601 18797 2635
rect 18797 2601 18831 2635
rect 18831 2601 18840 2635
rect 18788 2592 18840 2601
rect 8576 2524 8628 2576
rect 11612 2524 11664 2576
rect 16488 2524 16540 2576
rect 5816 2388 5868 2440
rect 6736 2431 6788 2440
rect 6736 2397 6745 2431
rect 6745 2397 6779 2431
rect 6779 2397 6788 2431
rect 6736 2388 6788 2397
rect 7104 2388 7156 2440
rect 7748 2388 7800 2440
rect 8116 2431 8168 2440
rect 8116 2397 8125 2431
rect 8125 2397 8159 2431
rect 8159 2397 8168 2431
rect 8116 2388 8168 2397
rect 9312 2431 9364 2440
rect 9312 2397 9321 2431
rect 9321 2397 9355 2431
rect 9355 2397 9364 2431
rect 9312 2388 9364 2397
rect 10600 2431 10652 2440
rect 10600 2397 10609 2431
rect 10609 2397 10643 2431
rect 10643 2397 10652 2431
rect 10600 2388 10652 2397
rect 10968 2388 11020 2440
rect 11704 2431 11756 2440
rect 11704 2397 11713 2431
rect 11713 2397 11747 2431
rect 11747 2397 11756 2431
rect 11704 2388 11756 2397
rect 12164 2431 12216 2440
rect 12164 2397 12173 2431
rect 12173 2397 12207 2431
rect 12207 2397 12216 2431
rect 12164 2388 12216 2397
rect 12256 2388 12308 2440
rect 13820 2431 13872 2440
rect 13820 2397 13829 2431
rect 13829 2397 13863 2431
rect 13863 2397 13872 2431
rect 13820 2388 13872 2397
rect 14464 2431 14516 2440
rect 14464 2397 14473 2431
rect 14473 2397 14507 2431
rect 14507 2397 14516 2431
rect 14464 2388 14516 2397
rect 15476 2388 15528 2440
rect 16672 2388 16724 2440
rect 17684 2431 17736 2440
rect 17684 2397 17693 2431
rect 17693 2397 17727 2431
rect 17727 2397 17736 2431
rect 17684 2388 17736 2397
rect 17960 2431 18012 2440
rect 17960 2397 17969 2431
rect 17969 2397 18003 2431
rect 18003 2397 18012 2431
rect 17960 2388 18012 2397
rect 18236 2431 18288 2440
rect 18236 2397 18245 2431
rect 18245 2397 18279 2431
rect 18279 2397 18288 2431
rect 18236 2388 18288 2397
rect 18512 2431 18564 2440
rect 18512 2397 18521 2431
rect 18521 2397 18555 2431
rect 18555 2397 18564 2431
rect 18512 2388 18564 2397
rect 18604 2431 18656 2440
rect 18604 2397 18613 2431
rect 18613 2397 18647 2431
rect 18647 2397 18656 2431
rect 18604 2388 18656 2397
rect 6460 2252 6512 2304
rect 9036 2252 9088 2304
rect 10324 2252 10376 2304
rect 12440 2252 12492 2304
rect 13544 2252 13596 2304
rect 14188 2252 14240 2304
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
<< metal2 >>
rect 5170 21706 5226 22401
rect 5814 21706 5870 22401
rect 6458 21706 6514 22401
rect 7102 21706 7158 22401
rect 7746 21706 7802 22401
rect 5170 21678 5304 21706
rect 5170 21601 5226 21678
rect 2350 20156 2658 20165
rect 2350 20154 2356 20156
rect 2412 20154 2436 20156
rect 2492 20154 2516 20156
rect 2572 20154 2596 20156
rect 2652 20154 2658 20156
rect 2412 20102 2414 20154
rect 2594 20102 2596 20154
rect 2350 20100 2356 20102
rect 2412 20100 2436 20102
rect 2492 20100 2516 20102
rect 2572 20100 2596 20102
rect 2652 20100 2658 20102
rect 2350 20091 2658 20100
rect 5276 20058 5304 21678
rect 5814 21678 5948 21706
rect 5814 21601 5870 21678
rect 5264 20052 5316 20058
rect 5264 19994 5316 20000
rect 5920 19854 5948 21678
rect 6458 21678 6776 21706
rect 6458 21601 6514 21678
rect 6748 19854 6776 21678
rect 7102 21678 7236 21706
rect 7102 21601 7158 21678
rect 7208 19854 7236 21678
rect 7576 21678 7802 21706
rect 4896 19848 4948 19854
rect 4896 19790 4948 19796
rect 5908 19848 5960 19854
rect 5908 19790 5960 19796
rect 6736 19848 6788 19854
rect 6736 19790 6788 19796
rect 7196 19848 7248 19854
rect 7196 19790 7248 19796
rect 3010 19612 3318 19621
rect 3010 19610 3016 19612
rect 3072 19610 3096 19612
rect 3152 19610 3176 19612
rect 3232 19610 3256 19612
rect 3312 19610 3318 19612
rect 3072 19558 3074 19610
rect 3254 19558 3256 19610
rect 3010 19556 3016 19558
rect 3072 19556 3096 19558
rect 3152 19556 3176 19558
rect 3232 19556 3256 19558
rect 3312 19556 3318 19558
rect 3010 19547 3318 19556
rect 4908 19514 4936 19790
rect 5724 19712 5776 19718
rect 5724 19654 5776 19660
rect 6552 19712 6604 19718
rect 6552 19654 6604 19660
rect 4896 19508 4948 19514
rect 4896 19450 4948 19456
rect 2872 19440 2924 19446
rect 2872 19382 2924 19388
rect 3976 19440 4028 19446
rect 3976 19382 4028 19388
rect 2688 19236 2740 19242
rect 2688 19178 2740 19184
rect 2350 19068 2658 19077
rect 2350 19066 2356 19068
rect 2412 19066 2436 19068
rect 2492 19066 2516 19068
rect 2572 19066 2596 19068
rect 2652 19066 2658 19068
rect 2412 19014 2414 19066
rect 2594 19014 2596 19066
rect 2350 19012 2356 19014
rect 2412 19012 2436 19014
rect 2492 19012 2516 19014
rect 2572 19012 2596 19014
rect 2652 19012 2658 19014
rect 2350 19003 2658 19012
rect 848 18760 900 18766
rect 848 18702 900 18708
rect 1676 18760 1728 18766
rect 1676 18702 1728 18708
rect 860 18601 888 18702
rect 846 18592 902 18601
rect 846 18527 902 18536
rect 1584 18080 1636 18086
rect 1584 18022 1636 18028
rect 1596 17882 1624 18022
rect 1584 17876 1636 17882
rect 1584 17818 1636 17824
rect 848 17672 900 17678
rect 846 17640 848 17649
rect 900 17640 902 17649
rect 846 17575 902 17584
rect 1216 17264 1268 17270
rect 1216 17206 1268 17212
rect 1228 17105 1256 17206
rect 1584 17196 1636 17202
rect 1584 17138 1636 17144
rect 1214 17096 1270 17105
rect 1214 17031 1270 17040
rect 1400 16992 1452 16998
rect 1400 16934 1452 16940
rect 1412 16425 1440 16934
rect 1596 16794 1624 17138
rect 1688 16794 1716 18702
rect 2320 18692 2372 18698
rect 2320 18634 2372 18640
rect 1768 18624 1820 18630
rect 1768 18566 1820 18572
rect 1780 18426 1808 18566
rect 2332 18426 2360 18634
rect 1768 18420 1820 18426
rect 1768 18362 1820 18368
rect 2320 18420 2372 18426
rect 2320 18362 2372 18368
rect 2596 18352 2648 18358
rect 2596 18294 2648 18300
rect 1952 18148 2004 18154
rect 1952 18090 2004 18096
rect 1584 16788 1636 16794
rect 1584 16730 1636 16736
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1688 16658 1716 16730
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 1584 16584 1636 16590
rect 1584 16526 1636 16532
rect 1398 16416 1454 16425
rect 1398 16351 1454 16360
rect 1596 16182 1624 16526
rect 1584 16176 1636 16182
rect 1584 16118 1636 16124
rect 848 16108 900 16114
rect 848 16050 900 16056
rect 860 15881 888 16050
rect 1768 15904 1820 15910
rect 846 15872 902 15881
rect 1768 15846 1820 15852
rect 846 15807 902 15816
rect 1400 15360 1452 15366
rect 1400 15302 1452 15308
rect 1412 15065 1440 15302
rect 1398 15056 1454 15065
rect 1398 14991 1454 15000
rect 1780 14958 1808 15846
rect 1860 15156 1912 15162
rect 1860 15098 1912 15104
rect 1676 14952 1728 14958
rect 1676 14894 1728 14900
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 1688 14482 1716 14894
rect 1676 14476 1728 14482
rect 1676 14418 1728 14424
rect 1780 14414 1808 14894
rect 1768 14408 1820 14414
rect 1030 14376 1086 14385
rect 1768 14350 1820 14356
rect 1030 14311 1086 14320
rect 1044 14006 1072 14311
rect 1676 14272 1728 14278
rect 1676 14214 1728 14220
rect 1768 14272 1820 14278
rect 1768 14214 1820 14220
rect 1688 14074 1716 14214
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 1032 14000 1084 14006
rect 1032 13942 1084 13948
rect 1492 13932 1544 13938
rect 1492 13874 1544 13880
rect 1504 13705 1532 13874
rect 1780 13802 1808 14214
rect 1768 13796 1820 13802
rect 1768 13738 1820 13744
rect 1490 13696 1546 13705
rect 1490 13631 1546 13640
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1214 13016 1270 13025
rect 1214 12951 1216 12960
rect 1268 12951 1270 12960
rect 1216 12922 1268 12928
rect 1596 12850 1624 13126
rect 1780 12850 1808 13738
rect 1872 13394 1900 15098
rect 1964 14550 1992 18090
rect 2608 18086 2636 18294
rect 2700 18290 2728 19178
rect 2688 18284 2740 18290
rect 2688 18226 2740 18232
rect 2780 18148 2832 18154
rect 2780 18090 2832 18096
rect 2228 18080 2280 18086
rect 2228 18022 2280 18028
rect 2596 18080 2648 18086
rect 2596 18022 2648 18028
rect 2240 17490 2268 18022
rect 2350 17980 2658 17989
rect 2350 17978 2356 17980
rect 2412 17978 2436 17980
rect 2492 17978 2516 17980
rect 2572 17978 2596 17980
rect 2652 17978 2658 17980
rect 2412 17926 2414 17978
rect 2594 17926 2596 17978
rect 2350 17924 2356 17926
rect 2412 17924 2436 17926
rect 2492 17924 2516 17926
rect 2572 17924 2596 17926
rect 2652 17924 2658 17926
rect 2350 17915 2658 17924
rect 2240 17462 2360 17490
rect 2332 17202 2360 17462
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 2320 17196 2372 17202
rect 2320 17138 2372 17144
rect 2044 16992 2096 16998
rect 2044 16934 2096 16940
rect 2056 16658 2084 16934
rect 2044 16652 2096 16658
rect 2044 16594 2096 16600
rect 2148 16114 2176 17138
rect 2228 17128 2280 17134
rect 2228 17070 2280 17076
rect 2240 16250 2268 17070
rect 2792 16998 2820 18090
rect 2780 16992 2832 16998
rect 2780 16934 2832 16940
rect 2350 16892 2658 16901
rect 2350 16890 2356 16892
rect 2412 16890 2436 16892
rect 2492 16890 2516 16892
rect 2572 16890 2596 16892
rect 2652 16890 2658 16892
rect 2412 16838 2414 16890
rect 2594 16838 2596 16890
rect 2350 16836 2356 16838
rect 2412 16836 2436 16838
rect 2492 16836 2516 16838
rect 2572 16836 2596 16838
rect 2652 16836 2658 16838
rect 2350 16827 2658 16836
rect 2792 16574 2820 16934
rect 2700 16546 2820 16574
rect 2228 16244 2280 16250
rect 2228 16186 2280 16192
rect 2700 16114 2728 16546
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 2792 16250 2820 16390
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 2884 16114 2912 19382
rect 3988 18970 4016 19382
rect 5736 19378 5764 19654
rect 6564 19514 6592 19654
rect 6552 19508 6604 19514
rect 6552 19450 6604 19456
rect 6644 19440 6696 19446
rect 6644 19382 6696 19388
rect 5724 19372 5776 19378
rect 5724 19314 5776 19320
rect 5908 19372 5960 19378
rect 5908 19314 5960 19320
rect 5078 19272 5134 19281
rect 5736 19242 5764 19314
rect 5078 19207 5134 19216
rect 5724 19236 5776 19242
rect 3976 18964 4028 18970
rect 3976 18906 4028 18912
rect 3976 18760 4028 18766
rect 3976 18702 4028 18708
rect 3424 18692 3476 18698
rect 3424 18634 3476 18640
rect 3010 18524 3318 18533
rect 3010 18522 3016 18524
rect 3072 18522 3096 18524
rect 3152 18522 3176 18524
rect 3232 18522 3256 18524
rect 3312 18522 3318 18524
rect 3072 18470 3074 18522
rect 3254 18470 3256 18522
rect 3010 18468 3016 18470
rect 3072 18468 3096 18470
rect 3152 18468 3176 18470
rect 3232 18468 3256 18470
rect 3312 18468 3318 18470
rect 3010 18459 3318 18468
rect 3436 18426 3464 18634
rect 3516 18624 3568 18630
rect 3516 18566 3568 18572
rect 3424 18420 3476 18426
rect 3424 18362 3476 18368
rect 2964 18284 3016 18290
rect 2964 18226 3016 18232
rect 3332 18284 3384 18290
rect 3332 18226 3384 18232
rect 2976 18086 3004 18226
rect 3344 18154 3372 18226
rect 3528 18222 3556 18566
rect 3988 18290 4016 18702
rect 4620 18692 4672 18698
rect 4620 18634 4672 18640
rect 4632 18426 4660 18634
rect 4620 18420 4672 18426
rect 4620 18362 4672 18368
rect 3976 18284 4028 18290
rect 3976 18226 4028 18232
rect 3516 18216 3568 18222
rect 3516 18158 3568 18164
rect 3332 18148 3384 18154
rect 3332 18090 3384 18096
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 3424 18080 3476 18086
rect 3424 18022 3476 18028
rect 3010 17436 3318 17445
rect 3010 17434 3016 17436
rect 3072 17434 3096 17436
rect 3152 17434 3176 17436
rect 3232 17434 3256 17436
rect 3312 17434 3318 17436
rect 3072 17382 3074 17434
rect 3254 17382 3256 17434
rect 3010 17380 3016 17382
rect 3072 17380 3096 17382
rect 3152 17380 3176 17382
rect 3232 17380 3256 17382
rect 3312 17380 3318 17382
rect 3010 17371 3318 17380
rect 3436 17082 3464 18022
rect 3528 17202 3556 18158
rect 3516 17196 3568 17202
rect 3516 17138 3568 17144
rect 3884 17128 3936 17134
rect 3436 17066 3556 17082
rect 3884 17070 3936 17076
rect 3436 17060 3568 17066
rect 3436 17054 3516 17060
rect 3516 17002 3568 17008
rect 3424 16448 3476 16454
rect 3424 16390 3476 16396
rect 3010 16348 3318 16357
rect 3010 16346 3016 16348
rect 3072 16346 3096 16348
rect 3152 16346 3176 16348
rect 3232 16346 3256 16348
rect 3312 16346 3318 16348
rect 3072 16294 3074 16346
rect 3254 16294 3256 16346
rect 3010 16292 3016 16294
rect 3072 16292 3096 16294
rect 3152 16292 3176 16294
rect 3232 16292 3256 16294
rect 3312 16292 3318 16294
rect 3010 16283 3318 16292
rect 3436 16182 3464 16390
rect 3424 16176 3476 16182
rect 3424 16118 3476 16124
rect 2136 16108 2188 16114
rect 2136 16050 2188 16056
rect 2688 16108 2740 16114
rect 2688 16050 2740 16056
rect 2872 16108 2924 16114
rect 2872 16050 2924 16056
rect 2700 15910 2728 16050
rect 2688 15904 2740 15910
rect 2688 15846 2740 15852
rect 2350 15804 2658 15813
rect 2350 15802 2356 15804
rect 2412 15802 2436 15804
rect 2492 15802 2516 15804
rect 2572 15802 2596 15804
rect 2652 15802 2658 15804
rect 2412 15750 2414 15802
rect 2594 15750 2596 15802
rect 2350 15748 2356 15750
rect 2412 15748 2436 15750
rect 2492 15748 2516 15750
rect 2572 15748 2596 15750
rect 2652 15748 2658 15750
rect 2350 15739 2658 15748
rect 2700 15366 2728 15846
rect 2136 15360 2188 15366
rect 2136 15302 2188 15308
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 1952 14544 2004 14550
rect 1952 14486 2004 14492
rect 2148 14414 2176 15302
rect 2884 15076 2912 16050
rect 3424 15496 3476 15502
rect 3424 15438 3476 15444
rect 3010 15260 3318 15269
rect 3010 15258 3016 15260
rect 3072 15258 3096 15260
rect 3152 15258 3176 15260
rect 3232 15258 3256 15260
rect 3312 15258 3318 15260
rect 3072 15206 3074 15258
rect 3254 15206 3256 15258
rect 3010 15204 3016 15206
rect 3072 15204 3096 15206
rect 3152 15204 3176 15206
rect 3232 15204 3256 15206
rect 3312 15204 3318 15206
rect 3010 15195 3318 15204
rect 3436 15162 3464 15438
rect 3424 15156 3476 15162
rect 3424 15098 3476 15104
rect 2964 15088 3016 15094
rect 2884 15048 2964 15076
rect 3528 15042 3556 17002
rect 3792 16992 3844 16998
rect 3792 16934 3844 16940
rect 3804 16658 3832 16934
rect 3896 16726 3924 17070
rect 3884 16720 3936 16726
rect 3884 16662 3936 16668
rect 3792 16652 3844 16658
rect 3792 16594 3844 16600
rect 4620 16584 4672 16590
rect 4620 16526 4672 16532
rect 4632 16454 4660 16526
rect 4896 16516 4948 16522
rect 4896 16458 4948 16464
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 4620 16448 4672 16454
rect 4620 16390 4672 16396
rect 4080 16182 4108 16390
rect 4068 16176 4120 16182
rect 4068 16118 4120 16124
rect 2964 15030 3016 15036
rect 2780 15020 2832 15026
rect 2780 14962 2832 14968
rect 3436 15014 3556 15042
rect 3700 15020 3752 15026
rect 2688 14952 2740 14958
rect 2688 14894 2740 14900
rect 2350 14716 2658 14725
rect 2350 14714 2356 14716
rect 2412 14714 2436 14716
rect 2492 14714 2516 14716
rect 2572 14714 2596 14716
rect 2652 14714 2658 14716
rect 2412 14662 2414 14714
rect 2594 14662 2596 14714
rect 2350 14660 2356 14662
rect 2412 14660 2436 14662
rect 2492 14660 2516 14662
rect 2572 14660 2596 14662
rect 2652 14660 2658 14662
rect 2350 14651 2658 14660
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2148 13938 2176 14350
rect 2700 14006 2728 14894
rect 2792 14618 2820 14962
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 3010 14172 3318 14181
rect 3010 14170 3016 14172
rect 3072 14170 3096 14172
rect 3152 14170 3176 14172
rect 3232 14170 3256 14172
rect 3312 14170 3318 14172
rect 3072 14118 3074 14170
rect 3254 14118 3256 14170
rect 3010 14116 3016 14118
rect 3072 14116 3096 14118
rect 3152 14116 3176 14118
rect 3232 14116 3256 14118
rect 3312 14116 3318 14118
rect 3010 14107 3318 14116
rect 2688 14000 2740 14006
rect 2688 13942 2740 13948
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 2148 13410 2176 13874
rect 3148 13728 3200 13734
rect 3148 13670 3200 13676
rect 2350 13628 2658 13637
rect 2350 13626 2356 13628
rect 2412 13626 2436 13628
rect 2492 13626 2516 13628
rect 2572 13626 2596 13628
rect 2652 13626 2658 13628
rect 2412 13574 2414 13626
rect 2594 13574 2596 13626
rect 2350 13572 2356 13574
rect 2412 13572 2436 13574
rect 2492 13572 2516 13574
rect 2572 13572 2596 13574
rect 2652 13572 2658 13574
rect 2350 13563 2658 13572
rect 1860 13388 1912 13394
rect 2148 13382 2268 13410
rect 1860 13330 1912 13336
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 1688 12345 1716 12786
rect 1674 12336 1730 12345
rect 1674 12271 1730 12280
rect 1780 11830 1808 12786
rect 1768 11824 1820 11830
rect 1768 11766 1820 11772
rect 1768 11688 1820 11694
rect 1872 11676 1900 13330
rect 2136 13252 2188 13258
rect 2136 13194 2188 13200
rect 2148 12986 2176 13194
rect 2136 12980 2188 12986
rect 2136 12922 2188 12928
rect 2136 11824 2188 11830
rect 2136 11766 2188 11772
rect 1820 11648 1900 11676
rect 1768 11630 1820 11636
rect 2148 11354 2176 11766
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2240 11150 2268 13382
rect 3160 13258 3188 13670
rect 3148 13252 3200 13258
rect 3148 13194 3200 13200
rect 2872 13184 2924 13190
rect 2872 13126 2924 13132
rect 2884 12850 2912 13126
rect 3010 13084 3318 13093
rect 3010 13082 3016 13084
rect 3072 13082 3096 13084
rect 3152 13082 3176 13084
rect 3232 13082 3256 13084
rect 3312 13082 3318 13084
rect 3072 13030 3074 13082
rect 3254 13030 3256 13082
rect 3010 13028 3016 13030
rect 3072 13028 3096 13030
rect 3152 13028 3176 13030
rect 3232 13028 3256 13030
rect 3312 13028 3318 13030
rect 3010 13019 3318 13028
rect 3436 12918 3464 15014
rect 3700 14962 3752 14968
rect 3792 15020 3844 15026
rect 3792 14962 3844 14968
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3516 14544 3568 14550
rect 3516 14486 3568 14492
rect 3528 14278 3556 14486
rect 3620 14346 3648 14758
rect 3712 14550 3740 14962
rect 3700 14544 3752 14550
rect 3700 14486 3752 14492
rect 3804 14482 3832 14962
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 4528 14952 4580 14958
rect 4528 14894 4580 14900
rect 4080 14618 4108 14894
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 4540 14414 4568 14894
rect 4344 14408 4396 14414
rect 4264 14368 4344 14396
rect 3608 14340 3660 14346
rect 3608 14282 3660 14288
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 3424 12912 3476 12918
rect 3424 12854 3476 12860
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 2350 12540 2658 12549
rect 2350 12538 2356 12540
rect 2412 12538 2436 12540
rect 2492 12538 2516 12540
rect 2572 12538 2596 12540
rect 2652 12538 2658 12540
rect 2412 12486 2414 12538
rect 2594 12486 2596 12538
rect 2350 12484 2356 12486
rect 2412 12484 2436 12486
rect 2492 12484 2516 12486
rect 2572 12484 2596 12486
rect 2652 12484 2658 12486
rect 2350 12475 2658 12484
rect 3010 11996 3318 12005
rect 3010 11994 3016 11996
rect 3072 11994 3096 11996
rect 3152 11994 3176 11996
rect 3232 11994 3256 11996
rect 3312 11994 3318 11996
rect 3072 11942 3074 11994
rect 3254 11942 3256 11994
rect 3010 11940 3016 11942
rect 3072 11940 3096 11942
rect 3152 11940 3176 11942
rect 3232 11940 3256 11942
rect 3312 11940 3318 11942
rect 3010 11931 3318 11940
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 2350 11452 2658 11461
rect 2350 11450 2356 11452
rect 2412 11450 2436 11452
rect 2492 11450 2516 11452
rect 2572 11450 2596 11452
rect 2652 11450 2658 11452
rect 2412 11398 2414 11450
rect 2594 11398 2596 11450
rect 2350 11396 2356 11398
rect 2412 11396 2436 11398
rect 2492 11396 2516 11398
rect 2572 11396 2596 11398
rect 2652 11396 2658 11398
rect 2350 11387 2658 11396
rect 3160 11286 3188 11494
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 1412 10985 1440 11086
rect 1584 11008 1636 11014
rect 1398 10976 1454 10985
rect 1584 10950 1636 10956
rect 1398 10911 1454 10920
rect 1596 10742 1624 10950
rect 2240 10826 2268 11086
rect 3528 11082 3556 14214
rect 4264 13938 4292 14368
rect 4344 14350 4396 14356
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4540 14278 4568 14350
rect 4528 14272 4580 14278
rect 4528 14214 4580 14220
rect 4632 13938 4660 16390
rect 4908 16250 4936 16458
rect 4896 16244 4948 16250
rect 4896 16186 4948 16192
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 4252 13932 4304 13938
rect 4252 13874 4304 13880
rect 4620 13932 4672 13938
rect 4620 13874 4672 13880
rect 3792 13524 3844 13530
rect 3792 13466 3844 13472
rect 3804 11665 3832 13466
rect 3896 13258 3924 13874
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 4080 13326 4108 13806
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4632 13394 4660 13670
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 3884 13252 3936 13258
rect 3884 13194 3936 13200
rect 3896 12102 3924 13194
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 3988 12850 4016 13126
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 4080 12782 4108 13262
rect 4068 12776 4120 12782
rect 4068 12718 4120 12724
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3896 11762 3924 12038
rect 4080 11762 4108 12718
rect 4436 12096 4488 12102
rect 4436 12038 4488 12044
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4172 11762 4200 11834
rect 4448 11762 4476 12038
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4816 11762 4844 11834
rect 5092 11830 5120 19207
rect 5724 19178 5776 19184
rect 5632 19168 5684 19174
rect 5632 19110 5684 19116
rect 5644 18698 5672 19110
rect 5632 18692 5684 18698
rect 5632 18634 5684 18640
rect 5736 16658 5764 19178
rect 5816 19168 5868 19174
rect 5816 19110 5868 19116
rect 5828 18426 5856 19110
rect 5816 18420 5868 18426
rect 5816 18362 5868 18368
rect 5920 18222 5948 19314
rect 6460 19168 6512 19174
rect 6460 19110 6512 19116
rect 6472 18698 6500 19110
rect 6552 18828 6604 18834
rect 6656 18816 6684 19382
rect 6736 19372 6788 19378
rect 6736 19314 6788 19320
rect 6604 18788 6684 18816
rect 6552 18770 6604 18776
rect 6460 18692 6512 18698
rect 6460 18634 6512 18640
rect 6000 18624 6052 18630
rect 6000 18566 6052 18572
rect 6012 18290 6040 18566
rect 6472 18358 6500 18634
rect 6460 18352 6512 18358
rect 6460 18294 6512 18300
rect 6000 18284 6052 18290
rect 6000 18226 6052 18232
rect 5908 18216 5960 18222
rect 5908 18158 5960 18164
rect 5920 18086 5948 18158
rect 5908 18080 5960 18086
rect 5908 18022 5960 18028
rect 6368 17672 6420 17678
rect 6368 17614 6420 17620
rect 6460 17672 6512 17678
rect 6460 17614 6512 17620
rect 6092 16992 6144 16998
rect 6092 16934 6144 16940
rect 5724 16652 5776 16658
rect 5724 16594 5776 16600
rect 6104 16590 6132 16934
rect 6380 16590 6408 17614
rect 6472 16794 6500 17614
rect 6564 17270 6592 18770
rect 6748 18714 6776 19314
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 7196 19168 7248 19174
rect 7196 19110 7248 19116
rect 6656 18686 6776 18714
rect 6552 17264 6604 17270
rect 6552 17206 6604 17212
rect 6460 16788 6512 16794
rect 6460 16730 6512 16736
rect 6564 16658 6592 17206
rect 6656 17202 6684 18686
rect 6840 18426 6868 19110
rect 7208 18698 7236 19110
rect 7196 18692 7248 18698
rect 7196 18634 7248 18640
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 6828 18420 6880 18426
rect 6828 18362 6880 18368
rect 7392 18290 7420 18566
rect 7576 18290 7604 21678
rect 7746 21601 7802 21678
rect 8390 21706 8446 22401
rect 9034 21706 9090 22401
rect 9678 21706 9734 22401
rect 10322 21706 10378 22401
rect 10966 21706 11022 22401
rect 8390 21678 8524 21706
rect 8390 21601 8446 21678
rect 8496 20058 8524 21678
rect 9034 21678 9168 21706
rect 9034 21601 9090 21678
rect 8484 20052 8536 20058
rect 8484 19994 8536 20000
rect 8668 19848 8720 19854
rect 8668 19790 8720 19796
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8404 18766 8432 19654
rect 8680 18970 8708 19790
rect 8760 19304 8812 19310
rect 8760 19246 8812 19252
rect 8772 18970 8800 19246
rect 8668 18964 8720 18970
rect 8668 18906 8720 18912
rect 8760 18964 8812 18970
rect 8760 18906 8812 18912
rect 9140 18834 9168 21678
rect 9678 21678 9812 21706
rect 9678 21601 9734 21678
rect 9784 20058 9812 21678
rect 10322 21678 10640 21706
rect 10322 21601 10378 21678
rect 9772 20052 9824 20058
rect 9772 19994 9824 20000
rect 10612 19854 10640 21678
rect 10888 21678 11022 21706
rect 10888 20058 10916 21678
rect 10966 21601 11022 21678
rect 11610 21706 11666 22401
rect 12254 21706 12310 22401
rect 12898 21706 12954 22401
rect 13542 21706 13598 22401
rect 14186 21706 14242 22401
rect 14830 21706 14886 22401
rect 16118 21706 16174 22401
rect 17498 21856 17554 21865
rect 17498 21791 17554 21800
rect 11610 21678 11744 21706
rect 11610 21601 11666 21678
rect 11716 20058 11744 21678
rect 12254 21678 12388 21706
rect 12254 21601 12310 21678
rect 10876 20052 10928 20058
rect 10876 19994 10928 20000
rect 11704 20052 11756 20058
rect 11704 19994 11756 20000
rect 9956 19848 10008 19854
rect 9956 19790 10008 19796
rect 10600 19848 10652 19854
rect 10600 19790 10652 19796
rect 11704 19848 11756 19854
rect 11704 19790 11756 19796
rect 9496 19780 9548 19786
rect 9496 19722 9548 19728
rect 9404 19712 9456 19718
rect 9404 19654 9456 19660
rect 9312 19440 9364 19446
rect 9312 19382 9364 19388
rect 9324 18970 9352 19382
rect 9312 18964 9364 18970
rect 9312 18906 9364 18912
rect 9128 18828 9180 18834
rect 9128 18770 9180 18776
rect 9416 18766 9444 19654
rect 9508 19514 9536 19722
rect 9496 19508 9548 19514
rect 9496 19450 9548 19456
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 8392 18760 8444 18766
rect 8392 18702 8444 18708
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7564 18284 7616 18290
rect 7564 18226 7616 18232
rect 6736 18216 6788 18222
rect 6736 18158 6788 18164
rect 6748 17814 6776 18158
rect 6736 17808 6788 17814
rect 6736 17750 6788 17756
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6092 16584 6144 16590
rect 6092 16526 6144 16532
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 6380 16454 6408 16526
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 6564 16046 6592 16594
rect 6656 16454 6684 17138
rect 6644 16448 6696 16454
rect 6644 16390 6696 16396
rect 6552 16040 6604 16046
rect 6552 15982 6604 15988
rect 5816 15904 5868 15910
rect 5816 15846 5868 15852
rect 5828 15502 5856 15846
rect 6564 15570 6592 15982
rect 6656 15706 6684 16390
rect 7392 16114 7420 18226
rect 7932 18080 7984 18086
rect 7932 18022 7984 18028
rect 7944 17270 7972 18022
rect 7932 17264 7984 17270
rect 7932 17206 7984 17212
rect 8300 16516 8352 16522
rect 8300 16458 8352 16464
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 7380 16108 7432 16114
rect 7380 16050 7432 16056
rect 6644 15700 6696 15706
rect 6644 15642 6696 15648
rect 6552 15564 6604 15570
rect 6552 15506 6604 15512
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 5724 15360 5776 15366
rect 5724 15302 5776 15308
rect 5736 15094 5764 15302
rect 5724 15088 5776 15094
rect 5724 15030 5776 15036
rect 5632 15020 5684 15026
rect 5632 14962 5684 14968
rect 5540 14816 5592 14822
rect 5540 14758 5592 14764
rect 5552 14346 5580 14758
rect 5644 14482 5672 14962
rect 5632 14476 5684 14482
rect 5632 14418 5684 14424
rect 5540 14340 5592 14346
rect 5540 14282 5592 14288
rect 5552 13870 5580 14282
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 5816 13864 5868 13870
rect 5816 13806 5868 13812
rect 5828 13530 5856 13806
rect 6000 13796 6052 13802
rect 6000 13738 6052 13744
rect 6012 13530 6040 13738
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 6656 13326 6684 15642
rect 6932 14822 6960 16050
rect 8116 16040 8168 16046
rect 8116 15982 8168 15988
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 7208 15162 7236 15302
rect 7300 15162 7328 15846
rect 8128 15706 8156 15982
rect 8116 15700 8168 15706
rect 8116 15642 8168 15648
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 7288 15156 7340 15162
rect 7288 15098 7340 15104
rect 7012 15088 7064 15094
rect 7012 15030 7064 15036
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 5356 12912 5408 12918
rect 5356 12854 5408 12860
rect 5080 11824 5132 11830
rect 5080 11766 5132 11772
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 4160 11756 4212 11762
rect 4160 11698 4212 11704
rect 4436 11756 4488 11762
rect 4436 11698 4488 11704
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 3790 11656 3846 11665
rect 4172 11642 4200 11698
rect 3790 11591 3846 11600
rect 4080 11614 4200 11642
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 3804 11286 3832 11591
rect 4080 11354 4108 11614
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 3792 11280 3844 11286
rect 3792 11222 3844 11228
rect 3884 11144 3936 11150
rect 3884 11086 3936 11092
rect 2780 11076 2832 11082
rect 2780 11018 2832 11024
rect 3516 11076 3568 11082
rect 3516 11018 3568 11024
rect 2148 10798 2268 10826
rect 1584 10736 1636 10742
rect 1584 10678 1636 10684
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 846 10160 902 10169
rect 846 10095 848 10104
rect 900 10095 902 10104
rect 848 10066 900 10072
rect 1412 9602 1440 10542
rect 2148 10062 2176 10798
rect 2228 10736 2280 10742
rect 2228 10678 2280 10684
rect 2240 10266 2268 10678
rect 2350 10364 2658 10373
rect 2350 10362 2356 10364
rect 2412 10362 2436 10364
rect 2492 10362 2516 10364
rect 2572 10362 2596 10364
rect 2652 10362 2658 10364
rect 2412 10310 2414 10362
rect 2594 10310 2596 10362
rect 2350 10308 2356 10310
rect 2412 10308 2436 10310
rect 2492 10308 2516 10310
rect 2572 10308 2596 10310
rect 2652 10308 2658 10310
rect 2350 10299 2658 10308
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 1412 9586 1532 9602
rect 848 9580 900 9586
rect 1412 9580 1544 9586
rect 1412 9574 1492 9580
rect 848 9522 900 9528
rect 1492 9522 1544 9528
rect 860 9489 888 9522
rect 846 9480 902 9489
rect 846 9415 902 9424
rect 848 9104 900 9110
rect 846 9072 848 9081
rect 900 9072 902 9081
rect 846 9007 902 9016
rect 2148 8974 2176 9998
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2350 9276 2658 9285
rect 2350 9274 2356 9276
rect 2412 9274 2436 9276
rect 2492 9274 2516 9276
rect 2572 9274 2596 9276
rect 2652 9274 2658 9276
rect 2412 9222 2414 9274
rect 2594 9222 2596 9274
rect 2350 9220 2356 9222
rect 2412 9220 2436 9222
rect 2492 9220 2516 9222
rect 2572 9220 2596 9222
rect 2652 9220 2658 9222
rect 2350 9211 2658 9220
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 1768 8288 1820 8294
rect 1306 8256 1362 8265
rect 1768 8230 1820 8236
rect 1306 8191 1362 8200
rect 1320 8090 1348 8191
rect 1308 8084 1360 8090
rect 1308 8026 1360 8032
rect 1780 7886 1808 8230
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 1872 7818 1900 8910
rect 2148 7886 2176 8910
rect 2700 8634 2728 9318
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2228 8560 2280 8566
rect 2228 8502 2280 8508
rect 2240 8090 2268 8502
rect 2350 8188 2658 8197
rect 2350 8186 2356 8188
rect 2412 8186 2436 8188
rect 2492 8186 2516 8188
rect 2572 8186 2596 8188
rect 2652 8186 2658 8188
rect 2412 8134 2414 8186
rect 2594 8134 2596 8186
rect 2350 8132 2356 8134
rect 2412 8132 2436 8134
rect 2492 8132 2516 8134
rect 2572 8132 2596 8134
rect 2652 8132 2658 8134
rect 2350 8123 2658 8132
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 2596 7880 2648 7886
rect 2648 7828 2728 7834
rect 2596 7822 2728 7828
rect 1860 7812 1912 7818
rect 2608 7806 2728 7822
rect 1860 7754 1912 7760
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 1306 7576 1362 7585
rect 1306 7511 1308 7520
rect 1360 7511 1362 7520
rect 1308 7482 1360 7488
rect 2516 7410 2544 7686
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2350 7100 2658 7109
rect 2350 7098 2356 7100
rect 2412 7098 2436 7100
rect 2492 7098 2516 7100
rect 2572 7098 2596 7100
rect 2652 7098 2658 7100
rect 2412 7046 2414 7098
rect 2594 7046 2596 7098
rect 2350 7044 2356 7046
rect 2412 7044 2436 7046
rect 2492 7044 2516 7046
rect 2572 7044 2596 7046
rect 2652 7044 2658 7046
rect 2350 7035 2658 7044
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 848 6316 900 6322
rect 848 6258 900 6264
rect 860 6089 888 6258
rect 846 6080 902 6089
rect 846 6015 902 6024
rect 1412 5778 1440 6734
rect 1676 6724 1728 6730
rect 1676 6666 1728 6672
rect 2412 6724 2464 6730
rect 2412 6666 2464 6672
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1412 5234 1440 5714
rect 1492 5568 1544 5574
rect 1490 5536 1492 5545
rect 1544 5536 1546 5545
rect 1490 5471 1546 5480
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 1596 4865 1624 6258
rect 1688 6186 1716 6666
rect 2424 6458 2452 6666
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2700 6322 2728 7806
rect 2792 6322 2820 11018
rect 3010 10908 3318 10917
rect 3010 10906 3016 10908
rect 3072 10906 3096 10908
rect 3152 10906 3176 10908
rect 3232 10906 3256 10908
rect 3312 10906 3318 10908
rect 3072 10854 3074 10906
rect 3254 10854 3256 10906
rect 3010 10852 3016 10854
rect 3072 10852 3096 10854
rect 3152 10852 3176 10854
rect 3232 10852 3256 10854
rect 3312 10852 3318 10854
rect 3010 10843 3318 10852
rect 3896 10810 3924 11086
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 3010 9820 3318 9829
rect 3010 9818 3016 9820
rect 3072 9818 3096 9820
rect 3152 9818 3176 9820
rect 3232 9818 3256 9820
rect 3312 9818 3318 9820
rect 3072 9766 3074 9818
rect 3254 9766 3256 9818
rect 3010 9764 3016 9766
rect 3072 9764 3096 9766
rect 3152 9764 3176 9766
rect 3232 9764 3256 9766
rect 3312 9764 3318 9766
rect 3010 9755 3318 9764
rect 4172 9654 4200 11494
rect 4724 11354 4752 11630
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 4908 11286 4936 11494
rect 4804 11280 4856 11286
rect 4804 11222 4856 11228
rect 4896 11280 4948 11286
rect 4896 11222 4948 11228
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4816 11098 4844 11222
rect 4896 11144 4948 11150
rect 4816 11092 4896 11098
rect 4816 11086 4948 11092
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 4160 9648 4212 9654
rect 4160 9590 4212 9596
rect 2884 9178 2912 9590
rect 4264 9382 4292 11086
rect 4816 11070 4936 11086
rect 4908 10810 4936 11070
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 4264 8498 4292 9318
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 2884 7546 2912 8366
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 4172 8022 4200 8298
rect 4160 8016 4212 8022
rect 4160 7958 4212 7964
rect 3884 7948 3936 7954
rect 3884 7890 3936 7896
rect 3976 7948 4028 7954
rect 3976 7890 4028 7896
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 1676 6180 1728 6186
rect 1676 6122 1728 6128
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 1768 5568 1820 5574
rect 1768 5510 1820 5516
rect 1780 5302 1808 5510
rect 1768 5296 1820 5302
rect 1768 5238 1820 5244
rect 1582 4856 1638 4865
rect 1582 4791 1638 4800
rect 1964 4690 1992 6054
rect 1952 4684 2004 4690
rect 1952 4626 2004 4632
rect 848 4616 900 4622
rect 848 4558 900 4564
rect 860 4321 888 4558
rect 846 4312 902 4321
rect 846 4247 902 4256
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 846 3632 902 3641
rect 846 3567 902 3576
rect 860 3534 888 3567
rect 848 3528 900 3534
rect 848 3470 900 3476
rect 1688 3194 1716 4082
rect 1964 4078 1992 4626
rect 2148 4622 2176 6258
rect 3436 6254 3464 6598
rect 3424 6248 3476 6254
rect 3424 6190 3476 6196
rect 2228 6180 2280 6186
rect 2228 6122 2280 6128
rect 2240 5710 2268 6122
rect 2350 6012 2658 6021
rect 2350 6010 2356 6012
rect 2412 6010 2436 6012
rect 2492 6010 2516 6012
rect 2572 6010 2596 6012
rect 2652 6010 2658 6012
rect 2412 5958 2414 6010
rect 2594 5958 2596 6010
rect 2350 5956 2356 5958
rect 2412 5956 2436 5958
rect 2492 5956 2516 5958
rect 2572 5956 2596 5958
rect 2652 5956 2658 5958
rect 2350 5947 2658 5956
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2332 5710 2360 5850
rect 2780 5840 2832 5846
rect 2780 5782 2832 5788
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 2240 5166 2268 5646
rect 2228 5160 2280 5166
rect 2228 5102 2280 5108
rect 2136 4616 2188 4622
rect 2136 4558 2188 4564
rect 2044 4548 2096 4554
rect 2044 4490 2096 4496
rect 2056 4146 2084 4490
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 1952 4072 2004 4078
rect 1952 4014 2004 4020
rect 2148 3738 2176 4558
rect 2240 4214 2268 5102
rect 2350 4924 2658 4933
rect 2350 4922 2356 4924
rect 2412 4922 2436 4924
rect 2492 4922 2516 4924
rect 2572 4922 2596 4924
rect 2652 4922 2658 4924
rect 2412 4870 2414 4922
rect 2594 4870 2596 4922
rect 2350 4868 2356 4870
rect 2412 4868 2436 4870
rect 2492 4868 2516 4870
rect 2572 4868 2596 4870
rect 2652 4868 2658 4870
rect 2350 4859 2658 4868
rect 2228 4208 2280 4214
rect 2228 4150 2280 4156
rect 2700 4078 2728 5714
rect 2792 5574 2820 5782
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 2780 5568 2832 5574
rect 2780 5510 2832 5516
rect 2792 5370 2820 5510
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 3528 5370 3556 5646
rect 3620 5642 3648 7822
rect 3896 7546 3924 7890
rect 3884 7540 3936 7546
rect 3884 7482 3936 7488
rect 3700 7404 3752 7410
rect 3700 7346 3752 7352
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3712 6866 3740 7346
rect 3792 7268 3844 7274
rect 3792 7210 3844 7216
rect 3700 6860 3752 6866
rect 3700 6802 3752 6808
rect 3804 6798 3832 7210
rect 3896 6882 3924 7346
rect 3988 7002 4016 7890
rect 4264 7410 4292 8298
rect 4540 7410 4568 10746
rect 5000 10606 5028 11698
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5264 11552 5316 11558
rect 5264 11494 5316 11500
rect 5092 11150 5120 11494
rect 5080 11144 5132 11150
rect 5080 11086 5132 11092
rect 5276 10742 5304 11494
rect 5368 11354 5396 12854
rect 6380 11762 6408 13262
rect 7024 12646 7052 15030
rect 8128 15026 8156 15642
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 8312 14414 8340 16458
rect 8404 16250 8432 18702
rect 9220 18284 9272 18290
rect 9220 18226 9272 18232
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8588 17270 8616 17478
rect 8576 17264 8628 17270
rect 8576 17206 8628 17212
rect 8680 16454 8708 17614
rect 9232 17338 9260 18226
rect 9220 17332 9272 17338
rect 9220 17274 9272 17280
rect 9600 17202 9628 19314
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9600 16658 9628 17138
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9220 16584 9272 16590
rect 9220 16526 9272 16532
rect 8668 16448 8720 16454
rect 8668 16390 8720 16396
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 8484 16176 8536 16182
rect 8484 16118 8536 16124
rect 8496 15706 8524 16118
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8680 15366 8708 16390
rect 9232 16250 9260 16526
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9508 16114 9536 16390
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 9692 15978 9720 18770
rect 9968 18426 9996 19790
rect 10508 19712 10560 19718
rect 10508 19654 10560 19660
rect 10232 19168 10284 19174
rect 10232 19110 10284 19116
rect 10244 18902 10272 19110
rect 10232 18896 10284 18902
rect 10232 18838 10284 18844
rect 10520 18698 10548 19654
rect 11716 19514 11744 19790
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 10968 19372 11020 19378
rect 10968 19314 11020 19320
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 10600 19304 10652 19310
rect 10600 19246 10652 19252
rect 10612 18970 10640 19246
rect 10980 18970 11008 19314
rect 10600 18964 10652 18970
rect 10600 18906 10652 18912
rect 10968 18964 11020 18970
rect 10968 18906 11020 18912
rect 10508 18692 10560 18698
rect 10508 18634 10560 18640
rect 9956 18420 10008 18426
rect 9956 18362 10008 18368
rect 10612 17678 10640 18906
rect 11152 18828 11204 18834
rect 11152 18770 11204 18776
rect 11164 18154 11192 18770
rect 11428 18624 11480 18630
rect 11428 18566 11480 18572
rect 11440 18358 11468 18566
rect 11428 18352 11480 18358
rect 11428 18294 11480 18300
rect 11152 18148 11204 18154
rect 11152 18090 11204 18096
rect 11164 17678 11192 18090
rect 11336 17740 11388 17746
rect 11336 17682 11388 17688
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 11152 17672 11204 17678
rect 11152 17614 11204 17620
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 9876 17270 9904 17478
rect 10796 17338 10824 17478
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 10888 17270 10916 17478
rect 9864 17264 9916 17270
rect 9864 17206 9916 17212
rect 10876 17264 10928 17270
rect 10876 17206 10928 17212
rect 11348 17134 11376 17682
rect 11440 17202 11468 18294
rect 11428 17196 11480 17202
rect 11428 17138 11480 17144
rect 11336 17128 11388 17134
rect 11336 17070 11388 17076
rect 10968 17060 11020 17066
rect 10968 17002 11020 17008
rect 10980 16658 11008 17002
rect 11440 16658 11468 17138
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 9680 15972 9732 15978
rect 9680 15914 9732 15920
rect 9312 15428 9364 15434
rect 9312 15370 9364 15376
rect 8668 15360 8720 15366
rect 8668 15302 8720 15308
rect 9324 15094 9352 15370
rect 11440 15094 11468 16594
rect 11532 15706 11560 19314
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 11704 18896 11756 18902
rect 11704 18838 11756 18844
rect 11716 18222 11744 18838
rect 11704 18216 11756 18222
rect 11704 18158 11756 18164
rect 11716 17202 11744 18158
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11520 15700 11572 15706
rect 11520 15642 11572 15648
rect 9312 15088 9364 15094
rect 9312 15030 9364 15036
rect 11428 15088 11480 15094
rect 11428 15030 11480 15036
rect 11440 14482 11468 15030
rect 11808 15026 11836 19110
rect 12164 18692 12216 18698
rect 12164 18634 12216 18640
rect 12176 18426 12204 18634
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 12360 18306 12388 21678
rect 12898 21678 13032 21706
rect 12898 21601 12954 21678
rect 13004 20058 13032 21678
rect 13542 21678 13768 21706
rect 13542 21601 13598 21678
rect 12992 20052 13044 20058
rect 12992 19994 13044 20000
rect 13740 19854 13768 21678
rect 14186 21678 14320 21706
rect 14186 21601 14242 21678
rect 14292 20058 14320 21678
rect 14830 21678 14964 21706
rect 14830 21601 14886 21678
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14936 19854 14964 21678
rect 16118 21678 16252 21706
rect 16118 21601 16174 21678
rect 16224 19854 16252 21678
rect 17512 20058 17540 21791
rect 17774 21176 17830 21185
rect 17774 21111 17830 21120
rect 17788 20058 17816 21111
rect 17958 20496 18014 20505
rect 17958 20431 18014 20440
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 17776 20052 17828 20058
rect 17776 19994 17828 20000
rect 13268 19848 13320 19854
rect 13268 19790 13320 19796
rect 13728 19848 13780 19854
rect 13728 19790 13780 19796
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 14924 19848 14976 19854
rect 14924 19790 14976 19796
rect 16212 19848 16264 19854
rect 16212 19790 16264 19796
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 12900 19712 12952 19718
rect 12900 19654 12952 19660
rect 12912 19378 12940 19654
rect 13280 19514 13308 19790
rect 14476 19514 14504 19790
rect 14924 19712 14976 19718
rect 14924 19654 14976 19660
rect 16396 19712 16448 19718
rect 16396 19654 16448 19660
rect 14936 19514 14964 19654
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 14464 19508 14516 19514
rect 14464 19450 14516 19456
rect 14924 19508 14976 19514
rect 14924 19450 14976 19456
rect 16408 19378 16436 19654
rect 17880 19514 17908 19790
rect 17868 19508 17920 19514
rect 17868 19450 17920 19456
rect 16948 19440 17000 19446
rect 16948 19382 17000 19388
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 13636 19372 13688 19378
rect 13636 19314 13688 19320
rect 15200 19372 15252 19378
rect 15200 19314 15252 19320
rect 16396 19372 16448 19378
rect 16396 19314 16448 19320
rect 12716 19168 12768 19174
rect 12716 19110 12768 19116
rect 12624 18828 12676 18834
rect 12624 18770 12676 18776
rect 12532 18308 12584 18314
rect 12360 18278 12532 18306
rect 12360 17882 12388 18278
rect 12532 18250 12584 18256
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 11900 17338 11928 17614
rect 11888 17332 11940 17338
rect 11888 17274 11940 17280
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 12268 16454 12296 17138
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 12452 16454 12480 17070
rect 12636 16794 12664 18770
rect 12728 18290 12756 19110
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 12912 18222 12940 19314
rect 13648 18970 13676 19314
rect 14832 19236 14884 19242
rect 14832 19178 14884 19184
rect 13636 18964 13688 18970
rect 13636 18906 13688 18912
rect 12992 18692 13044 18698
rect 12992 18634 13044 18640
rect 14648 18692 14700 18698
rect 14648 18634 14700 18640
rect 13004 18426 13032 18634
rect 14660 18426 14688 18634
rect 12992 18420 13044 18426
rect 12992 18362 13044 18368
rect 14648 18420 14700 18426
rect 14648 18362 14700 18368
rect 14844 18290 14872 19178
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 12716 18148 12768 18154
rect 12716 18090 12768 18096
rect 12728 16794 12756 18090
rect 15212 17626 15240 19314
rect 15292 19168 15344 19174
rect 15292 19110 15344 19116
rect 15304 18426 15332 19110
rect 16408 18766 16436 19314
rect 16672 19304 16724 19310
rect 16672 19246 16724 19252
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 15384 18692 15436 18698
rect 15384 18634 15436 18640
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15396 18154 15424 18634
rect 15660 18624 15712 18630
rect 15660 18566 15712 18572
rect 15672 18290 15700 18566
rect 15660 18284 15712 18290
rect 15660 18226 15712 18232
rect 15752 18216 15804 18222
rect 15752 18158 15804 18164
rect 15844 18216 15896 18222
rect 15844 18158 15896 18164
rect 15384 18148 15436 18154
rect 15384 18090 15436 18096
rect 15212 17610 15332 17626
rect 14832 17604 14884 17610
rect 15212 17604 15344 17610
rect 15212 17598 15292 17604
rect 14832 17546 14884 17552
rect 15292 17546 15344 17552
rect 14844 17338 14872 17546
rect 15200 17536 15252 17542
rect 15200 17478 15252 17484
rect 14832 17332 14884 17338
rect 14832 17274 14884 17280
rect 14924 17264 14976 17270
rect 14924 17206 14976 17212
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 13740 16794 13768 17138
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 12256 16448 12308 16454
rect 12256 16390 12308 16396
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12636 16250 12664 16730
rect 12728 16590 12756 16730
rect 14936 16590 14964 17206
rect 15212 17202 15240 17478
rect 15764 17338 15792 18158
rect 15856 17678 15884 18158
rect 16408 17746 16436 18702
rect 16488 18624 16540 18630
rect 16488 18566 16540 18572
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 16500 17678 16528 18566
rect 16684 18222 16712 19246
rect 16960 18970 16988 19382
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 16672 18216 16724 18222
rect 16672 18158 16724 18164
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16592 17785 16620 18022
rect 16578 17776 16634 17785
rect 16578 17711 16634 17720
rect 16592 17678 16620 17711
rect 16868 17678 16896 18702
rect 17684 18352 17736 18358
rect 17684 18294 17736 18300
rect 16948 18216 17000 18222
rect 16948 18158 17000 18164
rect 16960 17882 16988 18158
rect 17696 17882 17724 18294
rect 16948 17876 17000 17882
rect 16948 17818 17000 17824
rect 17684 17876 17736 17882
rect 17684 17818 17736 17824
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 15752 17332 15804 17338
rect 15752 17274 15804 17280
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15856 16658 15884 17614
rect 17776 17604 17828 17610
rect 17776 17546 17828 17552
rect 17788 17202 17816 17546
rect 17132 17196 17184 17202
rect 17132 17138 17184 17144
rect 17592 17196 17644 17202
rect 17592 17138 17644 17144
rect 17776 17196 17828 17202
rect 17776 17138 17828 17144
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 14924 16584 14976 16590
rect 14924 16526 14976 16532
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 12624 16244 12676 16250
rect 12624 16186 12676 16192
rect 12636 15502 12664 16186
rect 12728 15570 12756 16526
rect 14464 16448 14516 16454
rect 14464 16390 14516 16396
rect 14556 16448 14608 16454
rect 14556 16390 14608 16396
rect 13268 16176 13320 16182
rect 13268 16118 13320 16124
rect 13280 15706 13308 16118
rect 14188 16108 14240 16114
rect 14188 16050 14240 16056
rect 14096 16040 14148 16046
rect 14096 15982 14148 15988
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 13268 15700 13320 15706
rect 13268 15642 13320 15648
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 12624 15496 12676 15502
rect 12624 15438 12676 15444
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 13372 14550 13400 15846
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13360 14544 13412 14550
rect 13360 14486 13412 14492
rect 11428 14476 11480 14482
rect 11428 14418 11480 14424
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 10980 13258 11008 14350
rect 13372 13938 13400 14486
rect 13740 14414 13768 15438
rect 14108 15162 14136 15982
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 10968 13252 11020 13258
rect 10968 13194 11020 13200
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6380 11354 6408 11698
rect 10980 11558 11008 13194
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 13188 12782 13216 13126
rect 13372 12986 13400 13874
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 13924 12986 13952 13466
rect 14200 13326 14228 16050
rect 14372 15904 14424 15910
rect 14372 15846 14424 15852
rect 14384 15366 14412 15846
rect 14372 15360 14424 15366
rect 14372 15302 14424 15308
rect 14384 15026 14412 15302
rect 14476 15162 14504 16390
rect 14568 15502 14596 16390
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14936 15314 14964 16526
rect 15028 15706 15056 16526
rect 15856 16250 15884 16594
rect 17144 16454 17172 17138
rect 17604 17105 17632 17138
rect 17590 17096 17646 17105
rect 17590 17031 17646 17040
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 17328 16658 17356 16934
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 16212 16448 16264 16454
rect 16212 16390 16264 16396
rect 17132 16448 17184 16454
rect 17132 16390 17184 16396
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 15856 16130 15884 16186
rect 15856 16114 15976 16130
rect 15856 16108 15988 16114
rect 15856 16102 15936 16108
rect 15936 16050 15988 16056
rect 15016 15700 15068 15706
rect 15016 15642 15068 15648
rect 15948 15570 15976 16050
rect 16224 15570 16252 16390
rect 17144 15706 17172 16390
rect 17500 16176 17552 16182
rect 17500 16118 17552 16124
rect 17316 16040 17368 16046
rect 17316 15982 17368 15988
rect 17132 15700 17184 15706
rect 17132 15642 17184 15648
rect 15936 15564 15988 15570
rect 15936 15506 15988 15512
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 16764 15496 16816 15502
rect 16764 15438 16816 15444
rect 14936 15286 15148 15314
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 14372 15020 14424 15026
rect 14372 14962 14424 14968
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 14660 14414 14688 14554
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 14016 12986 14044 13262
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 13176 12776 13228 12782
rect 13176 12718 13228 12724
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 11900 12170 11928 12378
rect 13924 12306 13952 12922
rect 14292 12850 14320 14214
rect 14384 13870 14412 14350
rect 14464 14272 14516 14278
rect 14464 14214 14516 14220
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14476 13394 14504 14214
rect 15120 13818 15148 15286
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15660 14952 15712 14958
rect 15660 14894 15712 14900
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 15120 13790 15240 13818
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 14464 13388 14516 13394
rect 14464 13330 14516 13336
rect 15120 13258 15148 13466
rect 15108 13252 15160 13258
rect 15108 13194 15160 13200
rect 15212 12850 15240 13790
rect 15396 12866 15424 14214
rect 15488 12986 15516 14894
rect 15672 12986 15700 14894
rect 16028 14340 16080 14346
rect 16028 14282 16080 14288
rect 16040 13530 16068 14282
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16120 13864 16172 13870
rect 16120 13806 16172 13812
rect 16028 13524 16080 13530
rect 16028 13466 16080 13472
rect 16132 13326 16160 13806
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 15200 12844 15252 12850
rect 15396 12838 15608 12866
rect 15200 12786 15252 12792
rect 15108 12436 15160 12442
rect 15212 12434 15240 12786
rect 15160 12406 15240 12434
rect 15108 12378 15160 12384
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 11888 12164 11940 12170
rect 11888 12106 11940 12112
rect 12992 12164 13044 12170
rect 12992 12106 13044 12112
rect 14372 12164 14424 12170
rect 14372 12106 14424 12112
rect 15108 12164 15160 12170
rect 15108 12106 15160 12112
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 5552 10742 5580 11290
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5264 10736 5316 10742
rect 5264 10678 5316 10684
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 5828 10674 5856 11154
rect 6092 11076 6144 11082
rect 6092 11018 6144 11024
rect 6104 10810 6132 11018
rect 6092 10804 6144 10810
rect 6092 10746 6144 10752
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 4988 10600 5040 10606
rect 4988 10542 5040 10548
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5644 9042 5672 9318
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5828 8974 5856 10610
rect 6380 9586 6408 11290
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6840 11014 6868 11154
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6840 10810 6868 10950
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5828 8566 5856 8910
rect 5816 8560 5868 8566
rect 5816 8502 5868 8508
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4632 7478 4660 8434
rect 5828 7954 5856 8502
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4620 7472 4672 7478
rect 4620 7414 4672 7420
rect 4816 7410 4844 7686
rect 5552 7546 5580 7754
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 4528 7404 4580 7410
rect 4528 7346 4580 7352
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4264 7274 4292 7346
rect 4252 7268 4304 7274
rect 4252 7210 4304 7216
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 3896 6854 4016 6882
rect 4080 6866 4108 7142
rect 4264 7018 4292 7210
rect 4172 6990 4292 7018
rect 3988 6798 4016 6854
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 4066 6760 4122 6769
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3712 5846 3740 6258
rect 3700 5840 3752 5846
rect 3700 5782 3752 5788
rect 3608 5636 3660 5642
rect 3608 5578 3660 5584
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 2884 4826 2912 5170
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 3620 4690 3648 5170
rect 3608 4684 3660 4690
rect 3608 4626 3660 4632
rect 3712 4622 3740 5782
rect 3804 5710 3832 6734
rect 3896 5896 3924 6734
rect 3988 6458 4016 6734
rect 4172 6746 4200 6990
rect 5828 6866 5856 7890
rect 5920 7546 5948 9522
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 5920 7410 5948 7482
rect 6748 7426 6776 10542
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8116 9648 8168 9654
rect 8116 9590 8168 9596
rect 8128 8498 8156 9590
rect 8220 9058 8248 10066
rect 10612 9654 10640 11494
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 8220 9042 8340 9058
rect 8220 9036 8352 9042
rect 8220 9030 8300 9036
rect 8300 8978 8352 8984
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6840 7546 6868 7822
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 5908 7404 5960 7410
rect 6748 7398 6868 7426
rect 5908 7346 5960 7352
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 4122 6718 4200 6746
rect 4066 6695 4122 6704
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 3976 5908 4028 5914
rect 3896 5868 3976 5896
rect 3976 5850 4028 5856
rect 3988 5710 4016 5850
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 3804 5234 3832 5646
rect 3988 5302 4016 5646
rect 3976 5296 4028 5302
rect 3976 5238 4028 5244
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3804 4826 3832 5170
rect 4080 5098 4108 6695
rect 5920 5710 5948 7346
rect 6840 7274 6868 7398
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 6000 7268 6052 7274
rect 6000 7210 6052 7216
rect 6828 7268 6880 7274
rect 6828 7210 6880 7216
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 5816 5568 5868 5574
rect 5816 5510 5868 5516
rect 5828 5370 5856 5510
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 6012 5302 6040 7210
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6380 7002 6408 7142
rect 6368 6996 6420 7002
rect 6368 6938 6420 6944
rect 6840 5778 6868 7210
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 7116 6730 7144 7142
rect 7300 7002 7328 7346
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 7104 6724 7156 6730
rect 7104 6666 7156 6672
rect 7576 6254 7604 7278
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 6932 5574 6960 6190
rect 8024 5840 8076 5846
rect 8024 5782 8076 5788
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6000 5296 6052 5302
rect 6000 5238 6052 5244
rect 6932 5166 6960 5510
rect 7024 5234 7052 5646
rect 8036 5302 8064 5782
rect 8128 5710 8156 8434
rect 8312 7478 8340 8978
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 8588 8090 8616 8910
rect 9140 8634 9168 8910
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9324 8498 9352 8910
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 8312 6798 8340 7414
rect 8588 6798 8616 8026
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 9048 7478 9076 7686
rect 9036 7472 9088 7478
rect 9036 7414 9088 7420
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 9036 6792 9088 6798
rect 9036 6734 9088 6740
rect 8312 5914 8340 6734
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8588 5658 8616 6734
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 8864 5914 8892 6190
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 9048 5760 9076 6734
rect 9140 6322 9168 7822
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9508 6798 9536 7142
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9220 5772 9272 5778
rect 9048 5732 9220 5760
rect 8760 5704 8812 5710
rect 8588 5630 8708 5658
rect 8760 5646 8812 5652
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8024 5296 8076 5302
rect 8024 5238 8076 5244
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 7024 5114 7052 5170
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 5368 4622 5396 5102
rect 6932 4690 6960 5102
rect 7024 5086 7144 5114
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 4172 4282 4200 4422
rect 5368 4282 5396 4558
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 2350 3836 2658 3845
rect 2350 3834 2356 3836
rect 2412 3834 2436 3836
rect 2492 3834 2516 3836
rect 2572 3834 2596 3836
rect 2652 3834 2658 3836
rect 2412 3782 2414 3834
rect 2594 3782 2596 3834
rect 2350 3780 2356 3782
rect 2412 3780 2436 3782
rect 2492 3780 2516 3782
rect 2572 3780 2596 3782
rect 2652 3780 2658 3782
rect 2350 3771 2658 3780
rect 2136 3732 2188 3738
rect 2136 3674 2188 3680
rect 2700 3602 2728 4014
rect 2688 3596 2740 3602
rect 2688 3538 2740 3544
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 2700 3058 2728 3538
rect 3252 3534 3280 4082
rect 5552 3602 5580 4558
rect 6644 4480 6696 4486
rect 6696 4440 6776 4468
rect 6644 4422 6696 4428
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 3976 3392 4028 3398
rect 3976 3334 4028 3340
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 3988 3126 4016 3334
rect 3976 3120 4028 3126
rect 3976 3062 4028 3068
rect 5736 3058 5764 4082
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5828 3602 5856 3878
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 848 3052 900 3058
rect 848 2994 900 3000
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 860 2961 888 2994
rect 846 2952 902 2961
rect 6656 2922 6684 4082
rect 6748 3618 6776 4440
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6840 3738 6868 4082
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6932 3670 6960 4626
rect 7024 4554 7052 4966
rect 7012 4548 7064 4554
rect 7012 4490 7064 4496
rect 7116 4146 7144 5086
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7484 4146 7512 4966
rect 7668 4826 7696 5170
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 8116 4208 8168 4214
rect 8116 4150 8168 4156
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 6920 3664 6972 3670
rect 6748 3590 6868 3618
rect 6920 3606 6972 3612
rect 6840 3398 6868 3590
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 846 2887 902 2896
rect 6644 2916 6696 2922
rect 6644 2858 6696 2864
rect 6840 2854 6868 3334
rect 6932 3058 6960 3606
rect 7116 3466 7144 3878
rect 7300 3602 7328 4014
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 7104 3460 7156 3466
rect 7104 3402 7156 3408
rect 7012 3120 7064 3126
rect 7012 3062 7064 3068
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 6736 2848 6788 2854
rect 6736 2790 6788 2796
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 2350 2748 2658 2757
rect 2350 2746 2356 2748
rect 2412 2746 2436 2748
rect 2492 2746 2516 2748
rect 2572 2746 2596 2748
rect 2652 2746 2658 2748
rect 2412 2694 2414 2746
rect 2594 2694 2596 2746
rect 2350 2692 2356 2694
rect 2412 2692 2436 2694
rect 2492 2692 2516 2694
rect 2572 2692 2596 2694
rect 2652 2692 2658 2694
rect 2350 2683 2658 2692
rect 6748 2446 6776 2790
rect 6840 2650 6868 2790
rect 7024 2650 7052 3062
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 8128 2446 8156 4150
rect 8300 4004 8352 4010
rect 8300 3946 8352 3952
rect 8312 3534 8340 3946
rect 8392 3936 8444 3942
rect 8392 3878 8444 3884
rect 8404 3534 8432 3878
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8392 3528 8444 3534
rect 8444 3476 8524 3482
rect 8392 3470 8524 3476
rect 8404 3454 8524 3470
rect 8392 3120 8444 3126
rect 8392 3062 8444 3068
rect 8404 2650 8432 3062
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8496 2530 8524 3454
rect 8588 2582 8616 5510
rect 8680 4554 8708 5630
rect 8668 4548 8720 4554
rect 8668 4490 8720 4496
rect 8680 3602 8708 4490
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 8772 3194 8800 5646
rect 9048 5370 9076 5732
rect 9220 5714 9272 5720
rect 9324 5710 9352 6598
rect 9600 6458 9628 7278
rect 9692 7206 9720 8774
rect 9784 8498 9812 8774
rect 9876 8498 9904 8842
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 9600 5710 9628 6394
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 9588 5296 9640 5302
rect 9588 5238 9640 5244
rect 9600 4826 9628 5238
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8864 3534 8892 4082
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 9312 2848 9364 2854
rect 9312 2790 9364 2796
rect 8404 2502 8524 2530
rect 8576 2576 8628 2582
rect 8576 2518 8628 2524
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 5828 800 5856 2382
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 6472 800 6500 2246
rect 7116 800 7144 2382
rect 7760 800 7788 2382
rect 8404 800 8432 2502
rect 9324 2446 9352 2790
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 9048 800 9076 2246
rect 9692 800 9720 7142
rect 9784 6934 9812 7278
rect 9772 6928 9824 6934
rect 9772 6870 9824 6876
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9784 5710 9812 6258
rect 10968 5840 11020 5846
rect 10968 5782 11020 5788
rect 10980 5710 11008 5782
rect 11900 5778 11928 12106
rect 13004 11898 13032 12106
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 14384 11150 14412 12106
rect 15120 11898 15148 12106
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 15212 11762 15240 12406
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 15396 11286 15424 12038
rect 15384 11280 15436 11286
rect 15384 11222 15436 11228
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 11992 8838 12020 9522
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 12544 6390 12572 9590
rect 14200 9518 14228 10542
rect 15212 10266 15240 10542
rect 15200 10260 15252 10266
rect 15200 10202 15252 10208
rect 15396 9738 15424 11222
rect 15580 11150 15608 12838
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15672 11762 15700 12038
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15764 11558 15792 13262
rect 16500 12850 16528 14214
rect 16776 13938 16804 15438
rect 17328 15366 17356 15982
rect 17512 15706 17540 16118
rect 17500 15700 17552 15706
rect 17500 15642 17552 15648
rect 17604 15638 17632 17031
rect 17592 15632 17644 15638
rect 17592 15574 17644 15580
rect 17500 15496 17552 15502
rect 17500 15438 17552 15444
rect 17316 15360 17368 15366
rect 17316 15302 17368 15308
rect 17328 15094 17356 15302
rect 17316 15088 17368 15094
rect 17316 15030 17368 15036
rect 17040 15020 17092 15026
rect 17040 14962 17092 14968
rect 16948 14476 17000 14482
rect 17052 14464 17080 14962
rect 17316 14816 17368 14822
rect 17316 14758 17368 14764
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17328 14482 17356 14758
rect 17000 14436 17080 14464
rect 16948 14418 17000 14424
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16580 13932 16632 13938
rect 16580 13874 16632 13880
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 15844 11688 15896 11694
rect 15844 11630 15896 11636
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15764 11150 15792 11494
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15660 11076 15712 11082
rect 15660 11018 15712 11024
rect 15476 11008 15528 11014
rect 15476 10950 15528 10956
rect 15488 10062 15516 10950
rect 15672 10674 15700 11018
rect 15856 10810 15884 11630
rect 15936 11620 15988 11626
rect 15936 11562 15988 11568
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15856 10062 15884 10746
rect 15476 10056 15528 10062
rect 15476 9998 15528 10004
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 15396 9710 15516 9738
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14200 9382 14228 9454
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14200 8974 14228 9318
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 13740 7886 13768 8910
rect 14200 8498 14228 8910
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 14188 8492 14240 8498
rect 14108 8452 14188 8480
rect 14108 7954 14136 8452
rect 14188 8434 14240 8440
rect 15396 7954 15424 8774
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 15384 7948 15436 7954
rect 15384 7890 15436 7896
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 12532 6384 12584 6390
rect 12532 6326 12584 6332
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 13464 5710 13492 7822
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13740 6118 13768 7346
rect 14108 6866 14136 7890
rect 14648 7812 14700 7818
rect 14648 7754 14700 7760
rect 14660 7546 14688 7754
rect 14648 7540 14700 7546
rect 14648 7482 14700 7488
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15304 7410 15332 7482
rect 15396 7410 15424 7890
rect 15488 7410 15516 9710
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 15752 8424 15804 8430
rect 15752 8366 15804 8372
rect 15672 7970 15700 8366
rect 15764 8090 15792 8366
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 15672 7942 15792 7970
rect 15764 7750 15792 7942
rect 15948 7886 15976 11562
rect 16592 11370 16620 13874
rect 16868 13258 16896 14350
rect 17052 13734 17080 14436
rect 17316 14476 17368 14482
rect 17316 14418 17368 14424
rect 17420 14074 17448 14758
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17512 13870 17540 15438
rect 17788 15026 17816 17138
rect 17880 17066 17908 17614
rect 17868 17060 17920 17066
rect 17868 17002 17920 17008
rect 17880 15502 17908 17002
rect 17868 15496 17920 15502
rect 17868 15438 17920 15444
rect 17776 15020 17828 15026
rect 17776 14962 17828 14968
rect 17500 13864 17552 13870
rect 17500 13806 17552 13812
rect 17040 13728 17092 13734
rect 17040 13670 17092 13676
rect 17224 13728 17276 13734
rect 17224 13670 17276 13676
rect 17236 13394 17264 13670
rect 17224 13388 17276 13394
rect 17224 13330 17276 13336
rect 16856 13252 16908 13258
rect 16856 13194 16908 13200
rect 16868 12434 16896 13194
rect 16868 12406 16988 12434
rect 16960 11762 16988 12406
rect 17408 12164 17460 12170
rect 17408 12106 17460 12112
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 17224 11688 17276 11694
rect 17224 11630 17276 11636
rect 16500 11342 16620 11370
rect 17236 11354 17264 11630
rect 17224 11348 17276 11354
rect 16500 11286 16528 11342
rect 17224 11290 17276 11296
rect 17420 11286 17448 12106
rect 17592 12096 17644 12102
rect 17592 12038 17644 12044
rect 17500 11824 17552 11830
rect 17500 11766 17552 11772
rect 17512 11665 17540 11766
rect 17498 11656 17554 11665
rect 17498 11591 17554 11600
rect 16488 11280 16540 11286
rect 16488 11222 16540 11228
rect 17408 11280 17460 11286
rect 17408 11222 17460 11228
rect 17420 11150 17448 11222
rect 17512 11150 17540 11591
rect 17604 11150 17632 12038
rect 17788 11150 17816 14962
rect 17972 14890 18000 20431
rect 18236 19848 18288 19854
rect 18050 19816 18106 19825
rect 18236 19790 18288 19796
rect 18512 19848 18564 19854
rect 18512 19790 18564 19796
rect 18050 19751 18106 19760
rect 18064 19718 18092 19751
rect 18052 19712 18104 19718
rect 18052 19654 18104 19660
rect 18050 19136 18106 19145
rect 18050 19071 18106 19080
rect 18064 18970 18092 19071
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 18144 17536 18196 17542
rect 18144 17478 18196 17484
rect 18156 17202 18184 17478
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 18144 15904 18196 15910
rect 18144 15846 18196 15852
rect 18156 15026 18184 15846
rect 18248 15026 18276 19790
rect 18420 19168 18472 19174
rect 18420 19110 18472 19116
rect 18432 18766 18460 19110
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18340 18426 18368 18702
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18420 16992 18472 16998
rect 18420 16934 18472 16940
rect 18432 16590 18460 16934
rect 18420 16584 18472 16590
rect 18420 16526 18472 16532
rect 18524 16250 18552 19790
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18604 18624 18656 18630
rect 18604 18566 18656 18572
rect 18616 18290 18644 18566
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 18708 17270 18736 19314
rect 18786 18456 18842 18465
rect 18786 18391 18788 18400
rect 18840 18391 18842 18400
rect 18788 18362 18840 18368
rect 18788 17672 18840 17678
rect 18788 17614 18840 17620
rect 18696 17264 18748 17270
rect 18696 17206 18748 17212
rect 18708 16794 18736 17206
rect 18696 16788 18748 16794
rect 18696 16730 18748 16736
rect 18800 16425 18828 17614
rect 18786 16416 18842 16425
rect 18786 16351 18842 16360
rect 18512 16244 18564 16250
rect 18512 16186 18564 16192
rect 18788 16108 18840 16114
rect 18788 16050 18840 16056
rect 18800 15745 18828 16050
rect 18786 15736 18842 15745
rect 18786 15671 18842 15680
rect 18328 15496 18380 15502
rect 18328 15438 18380 15444
rect 18144 15020 18196 15026
rect 18144 14962 18196 14968
rect 18236 15020 18288 15026
rect 18236 14962 18288 14968
rect 17960 14884 18012 14890
rect 17960 14826 18012 14832
rect 18052 14340 18104 14346
rect 18052 14282 18104 14288
rect 18064 14074 18092 14282
rect 18248 14278 18276 14962
rect 18236 14272 18288 14278
rect 18236 14214 18288 14220
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 18340 12986 18368 15438
rect 18512 15428 18564 15434
rect 18512 15370 18564 15376
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 18432 13190 18460 13874
rect 18420 13184 18472 13190
rect 18420 13126 18472 13132
rect 18328 12980 18380 12986
rect 18328 12922 18380 12928
rect 18144 12844 18196 12850
rect 18144 12786 18196 12792
rect 18156 12238 18184 12786
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 17960 11824 18012 11830
rect 17960 11766 18012 11772
rect 17972 11354 18000 11766
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 18432 11150 18460 13126
rect 18524 12986 18552 15370
rect 18788 15360 18840 15366
rect 18788 15302 18840 15308
rect 18800 15065 18828 15302
rect 18786 15056 18842 15065
rect 18786 14991 18842 15000
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 18892 14385 18920 14962
rect 18878 14376 18934 14385
rect 18878 14311 18934 14320
rect 18788 14068 18840 14074
rect 18788 14010 18840 14016
rect 18604 13932 18656 13938
rect 18604 13874 18656 13880
rect 18616 13530 18644 13874
rect 18800 13705 18828 14010
rect 18786 13696 18842 13705
rect 18786 13631 18842 13640
rect 18604 13524 18656 13530
rect 18604 13466 18656 13472
rect 18786 13016 18842 13025
rect 18512 12980 18564 12986
rect 18786 12951 18842 12960
rect 18512 12922 18564 12928
rect 18800 12850 18828 12951
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 18786 12336 18842 12345
rect 18786 12271 18842 12280
rect 18800 12238 18828 12271
rect 18696 12232 18748 12238
rect 18696 12174 18748 12180
rect 18788 12232 18840 12238
rect 18788 12174 18840 12180
rect 18708 11898 18736 12174
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 17408 11144 17460 11150
rect 17408 11086 17460 11092
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17592 11144 17644 11150
rect 17776 11144 17828 11150
rect 17592 11086 17644 11092
rect 17696 11104 17776 11132
rect 16856 11008 16908 11014
rect 16856 10950 16908 10956
rect 16868 10130 16896 10950
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16592 9602 16620 9998
rect 16868 9994 16896 10066
rect 16856 9988 16908 9994
rect 16856 9930 16908 9936
rect 17408 9648 17460 9654
rect 16592 9574 16712 9602
rect 17408 9590 17460 9596
rect 16684 9518 16712 9574
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16028 8832 16080 8838
rect 16028 8774 16080 8780
rect 16040 7886 16068 8774
rect 15936 7880 15988 7886
rect 15936 7822 15988 7828
rect 16028 7880 16080 7886
rect 16028 7822 16080 7828
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15764 7478 15792 7686
rect 15752 7472 15804 7478
rect 15752 7414 15804 7420
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 14372 6792 14424 6798
rect 14648 6792 14700 6798
rect 14424 6740 14596 6746
rect 14372 6734 14596 6740
rect 14648 6734 14700 6740
rect 14384 6718 14596 6734
rect 14464 6656 14516 6662
rect 14464 6598 14516 6604
rect 14476 6458 14504 6598
rect 14568 6458 14596 6718
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14660 6322 14688 6734
rect 15304 6390 15332 7346
rect 15396 7206 15424 7346
rect 15844 7336 15896 7342
rect 15844 7278 15896 7284
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 15856 7002 15884 7278
rect 15844 6996 15896 7002
rect 15844 6938 15896 6944
rect 15568 6792 15620 6798
rect 15568 6734 15620 6740
rect 15292 6384 15344 6390
rect 15292 6326 15344 6332
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13740 5846 13768 6054
rect 14568 5914 14596 6258
rect 15016 6248 15068 6254
rect 15016 6190 15068 6196
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 13728 5840 13780 5846
rect 13728 5782 13780 5788
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 9784 4622 9812 5646
rect 13268 5636 13320 5642
rect 13268 5578 13320 5584
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 12072 5568 12124 5574
rect 12072 5510 12124 5516
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 10980 5302 11008 5510
rect 11244 5364 11296 5370
rect 11244 5306 11296 5312
rect 10968 5296 11020 5302
rect 10968 5238 11020 5244
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10704 4622 10732 4966
rect 11072 4826 11100 5102
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 9784 3618 9812 4558
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10704 3738 10732 4082
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 9784 3590 9904 3618
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9784 3194 9812 3402
rect 9876 3194 9904 3590
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9876 3058 9904 3130
rect 10704 3058 10732 3674
rect 10968 3120 11020 3126
rect 11020 3080 11100 3108
rect 10968 3062 11020 3068
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10600 2848 10652 2854
rect 10600 2790 10652 2796
rect 10612 2446 10640 2790
rect 11072 2650 11100 3080
rect 11164 2922 11192 4558
rect 11256 3058 11284 5306
rect 11428 5296 11480 5302
rect 11428 5238 11480 5244
rect 11440 4622 11468 5238
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 11336 4548 11388 4554
rect 11336 4490 11388 4496
rect 11348 4282 11376 4490
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 11440 3534 11468 4558
rect 11532 3602 11560 5102
rect 12084 4690 12112 5510
rect 12544 5302 12572 5510
rect 13280 5370 13308 5578
rect 13268 5364 13320 5370
rect 13268 5306 13320 5312
rect 12532 5296 12584 5302
rect 12532 5238 12584 5244
rect 12072 4684 12124 4690
rect 12072 4626 12124 4632
rect 12624 4480 12676 4486
rect 12624 4422 12676 4428
rect 12636 4146 12664 4422
rect 13464 4146 13492 5646
rect 13740 4622 13768 5782
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 14292 5302 14320 5646
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 14280 5296 14332 5302
rect 14280 5238 14332 5244
rect 14752 5234 14780 5510
rect 15028 5370 15056 6190
rect 15580 5778 15608 6734
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 15016 5364 15068 5370
rect 15016 5306 15068 5312
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 15948 5166 15976 7822
rect 16592 7750 16620 8910
rect 16684 8498 16712 9454
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16028 7404 16080 7410
rect 16028 7346 16080 7352
rect 16040 5846 16068 7346
rect 16592 6866 16620 7686
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16856 6724 16908 6730
rect 16856 6666 16908 6672
rect 16868 6458 16896 6666
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16960 6390 16988 9454
rect 17420 9178 17448 9590
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17408 8560 17460 8566
rect 17408 8502 17460 8508
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 17144 8090 17172 8366
rect 17420 8265 17448 8502
rect 17406 8256 17462 8265
rect 17406 8191 17462 8200
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 17420 7886 17448 8191
rect 17696 7886 17724 11104
rect 17776 11086 17828 11092
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 17972 9382 18000 10542
rect 18340 10266 18368 10610
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18432 10062 18460 11086
rect 18800 10985 18828 11086
rect 18786 10976 18842 10985
rect 18786 10911 18842 10920
rect 18604 10464 18656 10470
rect 18604 10406 18656 10412
rect 18788 10464 18840 10470
rect 18788 10406 18840 10412
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 17960 9376 18012 9382
rect 17960 9318 18012 9324
rect 18328 9376 18380 9382
rect 18328 9318 18380 9324
rect 18340 8974 18368 9318
rect 18616 8974 18644 10406
rect 18800 10305 18828 10406
rect 18786 10296 18842 10305
rect 18786 10231 18842 10240
rect 18786 9616 18842 9625
rect 18786 9551 18842 9560
rect 18800 9178 18828 9551
rect 18788 9172 18840 9178
rect 18788 9114 18840 9120
rect 18328 8968 18380 8974
rect 18604 8968 18656 8974
rect 18328 8910 18380 8916
rect 18510 8936 18566 8945
rect 18604 8910 18656 8916
rect 18510 8871 18566 8880
rect 18524 8838 18552 8871
rect 18512 8832 18564 8838
rect 18512 8774 18564 8780
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 18144 8288 18196 8294
rect 18144 8230 18196 8236
rect 18156 7886 18184 8230
rect 18248 8090 18276 8434
rect 18236 8084 18288 8090
rect 18236 8026 18288 8032
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 17696 7546 17724 7822
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17408 7472 17460 7478
rect 17408 7414 17460 7420
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 16580 6384 16632 6390
rect 16580 6326 16632 6332
rect 16948 6384 17000 6390
rect 16948 6326 17000 6332
rect 16592 5914 16620 6326
rect 17236 6322 17264 6802
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 16580 5908 16632 5914
rect 16580 5850 16632 5856
rect 16028 5840 16080 5846
rect 16028 5782 16080 5788
rect 15936 5160 15988 5166
rect 15936 5102 15988 5108
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 11900 3738 11928 4082
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 11992 3618 12020 4014
rect 12900 4004 12952 4010
rect 12900 3946 12952 3952
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 12268 3738 12296 3878
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 11900 3590 12020 3618
rect 11428 3528 11480 3534
rect 11428 3470 11480 3476
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11440 2922 11468 3470
rect 11532 3058 11560 3538
rect 11900 3534 11928 3590
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 11152 2916 11204 2922
rect 11152 2858 11204 2864
rect 11428 2916 11480 2922
rect 11428 2858 11480 2864
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11612 2576 11664 2582
rect 11612 2518 11664 2524
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 10336 800 10364 2246
rect 10980 800 11008 2382
rect 11624 800 11652 2518
rect 11716 2446 11744 3130
rect 11900 2990 11928 3470
rect 12072 3120 12124 3126
rect 12532 3120 12584 3126
rect 12124 3080 12296 3108
rect 12072 3062 12124 3068
rect 11888 2984 11940 2990
rect 11888 2926 11940 2932
rect 12268 2854 12296 3080
rect 12532 3062 12584 3068
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12164 2848 12216 2854
rect 12164 2790 12216 2796
rect 12256 2848 12308 2854
rect 12256 2790 12308 2796
rect 12176 2446 12204 2790
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 12268 800 12296 2382
rect 12452 2310 12480 2926
rect 12544 2650 12572 3062
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12912 800 12940 3946
rect 13004 3738 13032 4082
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 13464 3466 13492 3878
rect 13740 3602 13768 4558
rect 15396 4554 15424 4966
rect 15948 4622 15976 5102
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 15384 4548 15436 4554
rect 15384 4490 15436 4496
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 14384 3466 14412 3878
rect 13452 3460 13504 3466
rect 13452 3402 13504 3408
rect 14372 3460 14424 3466
rect 14372 3402 14424 3408
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13740 3058 13768 3334
rect 15212 3194 15240 4082
rect 15844 4072 15896 4078
rect 15844 4014 15896 4020
rect 15856 3738 15884 4014
rect 15936 4004 15988 4010
rect 15936 3946 15988 3952
rect 15948 3738 15976 3946
rect 15844 3732 15896 3738
rect 15844 3674 15896 3680
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 15844 3460 15896 3466
rect 15844 3402 15896 3408
rect 15856 3194 15884 3402
rect 15200 3188 15252 3194
rect 15200 3130 15252 3136
rect 15844 3188 15896 3194
rect 15844 3130 15896 3136
rect 15476 3120 15528 3126
rect 15476 3062 15528 3068
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 14464 2848 14516 2854
rect 14464 2790 14516 2796
rect 13832 2446 13860 2790
rect 14476 2446 14504 2790
rect 15488 2650 15516 3062
rect 16040 2990 16068 5782
rect 17132 5636 17184 5642
rect 17132 5578 17184 5584
rect 16488 5568 16540 5574
rect 16488 5510 16540 5516
rect 16396 4820 16448 4826
rect 16396 4762 16448 4768
rect 16408 4146 16436 4762
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16028 2984 16080 2990
rect 16028 2926 16080 2932
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 16500 2582 16528 5510
rect 17144 5370 17172 5578
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 17236 5302 17264 6258
rect 17316 6112 17368 6118
rect 17316 6054 17368 6060
rect 17224 5296 17276 5302
rect 17224 5238 17276 5244
rect 17132 5228 17184 5234
rect 17132 5170 17184 5176
rect 17144 5030 17172 5170
rect 17236 5166 17264 5238
rect 17224 5160 17276 5166
rect 17224 5102 17276 5108
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 16592 3534 16620 4422
rect 17040 4072 17092 4078
rect 17040 4014 17092 4020
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16592 2854 16620 3470
rect 16672 3460 16724 3466
rect 16672 3402 16724 3408
rect 16684 2922 16712 3402
rect 17052 3398 17080 4014
rect 17236 3466 17264 5102
rect 17328 5098 17356 6054
rect 17316 5092 17368 5098
rect 17316 5034 17368 5040
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17328 3738 17356 4014
rect 17316 3732 17368 3738
rect 17316 3674 17368 3680
rect 17224 3460 17276 3466
rect 17224 3402 17276 3408
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 16960 2990 16988 3130
rect 17052 3126 17080 3334
rect 17040 3120 17092 3126
rect 17040 3062 17092 3068
rect 17224 3120 17276 3126
rect 17224 3062 17276 3068
rect 16948 2984 17000 2990
rect 16948 2926 17000 2932
rect 16672 2916 16724 2922
rect 16672 2858 16724 2864
rect 16580 2848 16632 2854
rect 16580 2790 16632 2796
rect 16488 2576 16540 2582
rect 16488 2518 16540 2524
rect 16684 2446 16712 2858
rect 17236 2650 17264 3062
rect 17420 2650 17448 7414
rect 17500 6180 17552 6186
rect 17500 6122 17552 6128
rect 17512 5234 17540 6122
rect 17696 5234 17724 7482
rect 18064 6458 18092 7822
rect 18156 7410 18184 7822
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 18328 7404 18380 7410
rect 18328 7346 18380 7352
rect 18340 7002 18368 7346
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 18328 6996 18380 7002
rect 18328 6938 18380 6944
rect 18052 6452 18104 6458
rect 18052 6394 18104 6400
rect 17868 6316 17920 6322
rect 17868 6258 17920 6264
rect 17880 5778 17908 6258
rect 17868 5772 17920 5778
rect 17868 5714 17920 5720
rect 17500 5228 17552 5234
rect 17500 5170 17552 5176
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17590 4856 17646 4865
rect 17590 4791 17646 4800
rect 17696 4808 17724 5170
rect 17880 5030 17908 5714
rect 18144 5636 18196 5642
rect 18144 5578 18196 5584
rect 18156 5370 18184 5578
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 18524 5234 18552 7142
rect 18616 7002 18644 7822
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18800 7585 18828 7686
rect 18786 7576 18842 7585
rect 18786 7511 18842 7520
rect 18788 7200 18840 7206
rect 18788 7142 18840 7148
rect 18604 6996 18656 7002
rect 18604 6938 18656 6944
rect 18800 6905 18828 7142
rect 18786 6896 18842 6905
rect 18786 6831 18842 6840
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18616 6322 18644 6734
rect 18604 6316 18656 6322
rect 18604 6258 18656 6264
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18616 5914 18644 6258
rect 18800 6225 18828 6258
rect 18786 6216 18842 6225
rect 18786 6151 18842 6160
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18786 5536 18842 5545
rect 18786 5471 18842 5480
rect 18800 5370 18828 5471
rect 18788 5364 18840 5370
rect 18788 5306 18840 5312
rect 18512 5228 18564 5234
rect 18512 5170 18564 5176
rect 18144 5092 18196 5098
rect 18144 5034 18196 5040
rect 17868 5024 17920 5030
rect 17868 4966 17920 4972
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 17500 3936 17552 3942
rect 17604 3890 17632 4791
rect 17696 4780 17908 4808
rect 17776 4616 17828 4622
rect 17776 4558 17828 4564
rect 17684 4480 17736 4486
rect 17684 4422 17736 4428
rect 17552 3884 17632 3890
rect 17500 3878 17632 3884
rect 17512 3862 17632 3878
rect 17604 3534 17632 3862
rect 17696 3534 17724 4422
rect 17788 3602 17816 4558
rect 17880 3670 17908 4780
rect 17868 3664 17920 3670
rect 17868 3606 17920 3612
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 17684 3528 17736 3534
rect 17684 3470 17736 3476
rect 17788 2650 17816 3538
rect 17880 3534 17908 3606
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 18064 2650 18092 4966
rect 17224 2644 17276 2650
rect 17224 2586 17276 2592
rect 17408 2644 17460 2650
rect 17408 2586 17460 2592
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 14464 2440 14516 2446
rect 14464 2382 14516 2388
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 16672 2440 16724 2446
rect 16672 2382 16724 2388
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 17960 2440 18012 2446
rect 17960 2382 18012 2388
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 13556 800 13584 2246
rect 14200 800 14228 2246
rect 15488 800 15516 2382
rect 17696 1465 17724 2382
rect 17682 1456 17738 1465
rect 17682 1391 17738 1400
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 17972 785 18000 2382
rect 18156 2145 18184 5034
rect 18236 4616 18288 4622
rect 18236 4558 18288 4564
rect 18328 4616 18380 4622
rect 18328 4558 18380 4564
rect 18248 3602 18276 4558
rect 18340 3738 18368 4558
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 18800 4185 18828 4422
rect 18786 4176 18842 4185
rect 18420 4140 18472 4146
rect 18786 4111 18842 4120
rect 18420 4082 18472 4088
rect 18432 3738 18460 4082
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18328 3732 18380 3738
rect 18328 3674 18380 3680
rect 18420 3732 18472 3738
rect 18420 3674 18472 3680
rect 18800 3602 18828 3878
rect 18236 3596 18288 3602
rect 18236 3538 18288 3544
rect 18788 3596 18840 3602
rect 18788 3538 18840 3544
rect 18786 3496 18842 3505
rect 18786 3431 18842 3440
rect 18604 2848 18656 2854
rect 18510 2816 18566 2825
rect 18604 2790 18656 2796
rect 18510 2751 18566 2760
rect 18524 2446 18552 2751
rect 18616 2446 18644 2790
rect 18800 2650 18828 3431
rect 18788 2644 18840 2650
rect 18788 2586 18840 2592
rect 18236 2440 18288 2446
rect 18236 2382 18288 2388
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18604 2440 18656 2446
rect 18604 2382 18656 2388
rect 18142 2136 18198 2145
rect 18142 2071 18198 2080
rect 17958 776 18014 785
rect 17958 711 18014 720
rect 18050 0 18106 800
rect 18248 105 18276 2382
rect 18234 96 18290 105
rect 18234 31 18290 40
<< via2 >>
rect 2356 20154 2412 20156
rect 2436 20154 2492 20156
rect 2516 20154 2572 20156
rect 2596 20154 2652 20156
rect 2356 20102 2402 20154
rect 2402 20102 2412 20154
rect 2436 20102 2466 20154
rect 2466 20102 2478 20154
rect 2478 20102 2492 20154
rect 2516 20102 2530 20154
rect 2530 20102 2542 20154
rect 2542 20102 2572 20154
rect 2596 20102 2606 20154
rect 2606 20102 2652 20154
rect 2356 20100 2412 20102
rect 2436 20100 2492 20102
rect 2516 20100 2572 20102
rect 2596 20100 2652 20102
rect 3016 19610 3072 19612
rect 3096 19610 3152 19612
rect 3176 19610 3232 19612
rect 3256 19610 3312 19612
rect 3016 19558 3062 19610
rect 3062 19558 3072 19610
rect 3096 19558 3126 19610
rect 3126 19558 3138 19610
rect 3138 19558 3152 19610
rect 3176 19558 3190 19610
rect 3190 19558 3202 19610
rect 3202 19558 3232 19610
rect 3256 19558 3266 19610
rect 3266 19558 3312 19610
rect 3016 19556 3072 19558
rect 3096 19556 3152 19558
rect 3176 19556 3232 19558
rect 3256 19556 3312 19558
rect 2356 19066 2412 19068
rect 2436 19066 2492 19068
rect 2516 19066 2572 19068
rect 2596 19066 2652 19068
rect 2356 19014 2402 19066
rect 2402 19014 2412 19066
rect 2436 19014 2466 19066
rect 2466 19014 2478 19066
rect 2478 19014 2492 19066
rect 2516 19014 2530 19066
rect 2530 19014 2542 19066
rect 2542 19014 2572 19066
rect 2596 19014 2606 19066
rect 2606 19014 2652 19066
rect 2356 19012 2412 19014
rect 2436 19012 2492 19014
rect 2516 19012 2572 19014
rect 2596 19012 2652 19014
rect 846 18536 902 18592
rect 846 17620 848 17640
rect 848 17620 900 17640
rect 900 17620 902 17640
rect 846 17584 902 17620
rect 1214 17040 1270 17096
rect 1398 16360 1454 16416
rect 846 15816 902 15872
rect 1398 15000 1454 15056
rect 1030 14320 1086 14376
rect 1490 13640 1546 13696
rect 1214 12980 1270 13016
rect 1214 12960 1216 12980
rect 1216 12960 1268 12980
rect 1268 12960 1270 12980
rect 2356 17978 2412 17980
rect 2436 17978 2492 17980
rect 2516 17978 2572 17980
rect 2596 17978 2652 17980
rect 2356 17926 2402 17978
rect 2402 17926 2412 17978
rect 2436 17926 2466 17978
rect 2466 17926 2478 17978
rect 2478 17926 2492 17978
rect 2516 17926 2530 17978
rect 2530 17926 2542 17978
rect 2542 17926 2572 17978
rect 2596 17926 2606 17978
rect 2606 17926 2652 17978
rect 2356 17924 2412 17926
rect 2436 17924 2492 17926
rect 2516 17924 2572 17926
rect 2596 17924 2652 17926
rect 2356 16890 2412 16892
rect 2436 16890 2492 16892
rect 2516 16890 2572 16892
rect 2596 16890 2652 16892
rect 2356 16838 2402 16890
rect 2402 16838 2412 16890
rect 2436 16838 2466 16890
rect 2466 16838 2478 16890
rect 2478 16838 2492 16890
rect 2516 16838 2530 16890
rect 2530 16838 2542 16890
rect 2542 16838 2572 16890
rect 2596 16838 2606 16890
rect 2606 16838 2652 16890
rect 2356 16836 2412 16838
rect 2436 16836 2492 16838
rect 2516 16836 2572 16838
rect 2596 16836 2652 16838
rect 5078 19216 5134 19272
rect 3016 18522 3072 18524
rect 3096 18522 3152 18524
rect 3176 18522 3232 18524
rect 3256 18522 3312 18524
rect 3016 18470 3062 18522
rect 3062 18470 3072 18522
rect 3096 18470 3126 18522
rect 3126 18470 3138 18522
rect 3138 18470 3152 18522
rect 3176 18470 3190 18522
rect 3190 18470 3202 18522
rect 3202 18470 3232 18522
rect 3256 18470 3266 18522
rect 3266 18470 3312 18522
rect 3016 18468 3072 18470
rect 3096 18468 3152 18470
rect 3176 18468 3232 18470
rect 3256 18468 3312 18470
rect 3016 17434 3072 17436
rect 3096 17434 3152 17436
rect 3176 17434 3232 17436
rect 3256 17434 3312 17436
rect 3016 17382 3062 17434
rect 3062 17382 3072 17434
rect 3096 17382 3126 17434
rect 3126 17382 3138 17434
rect 3138 17382 3152 17434
rect 3176 17382 3190 17434
rect 3190 17382 3202 17434
rect 3202 17382 3232 17434
rect 3256 17382 3266 17434
rect 3266 17382 3312 17434
rect 3016 17380 3072 17382
rect 3096 17380 3152 17382
rect 3176 17380 3232 17382
rect 3256 17380 3312 17382
rect 3016 16346 3072 16348
rect 3096 16346 3152 16348
rect 3176 16346 3232 16348
rect 3256 16346 3312 16348
rect 3016 16294 3062 16346
rect 3062 16294 3072 16346
rect 3096 16294 3126 16346
rect 3126 16294 3138 16346
rect 3138 16294 3152 16346
rect 3176 16294 3190 16346
rect 3190 16294 3202 16346
rect 3202 16294 3232 16346
rect 3256 16294 3266 16346
rect 3266 16294 3312 16346
rect 3016 16292 3072 16294
rect 3096 16292 3152 16294
rect 3176 16292 3232 16294
rect 3256 16292 3312 16294
rect 2356 15802 2412 15804
rect 2436 15802 2492 15804
rect 2516 15802 2572 15804
rect 2596 15802 2652 15804
rect 2356 15750 2402 15802
rect 2402 15750 2412 15802
rect 2436 15750 2466 15802
rect 2466 15750 2478 15802
rect 2478 15750 2492 15802
rect 2516 15750 2530 15802
rect 2530 15750 2542 15802
rect 2542 15750 2572 15802
rect 2596 15750 2606 15802
rect 2606 15750 2652 15802
rect 2356 15748 2412 15750
rect 2436 15748 2492 15750
rect 2516 15748 2572 15750
rect 2596 15748 2652 15750
rect 3016 15258 3072 15260
rect 3096 15258 3152 15260
rect 3176 15258 3232 15260
rect 3256 15258 3312 15260
rect 3016 15206 3062 15258
rect 3062 15206 3072 15258
rect 3096 15206 3126 15258
rect 3126 15206 3138 15258
rect 3138 15206 3152 15258
rect 3176 15206 3190 15258
rect 3190 15206 3202 15258
rect 3202 15206 3232 15258
rect 3256 15206 3266 15258
rect 3266 15206 3312 15258
rect 3016 15204 3072 15206
rect 3096 15204 3152 15206
rect 3176 15204 3232 15206
rect 3256 15204 3312 15206
rect 2356 14714 2412 14716
rect 2436 14714 2492 14716
rect 2516 14714 2572 14716
rect 2596 14714 2652 14716
rect 2356 14662 2402 14714
rect 2402 14662 2412 14714
rect 2436 14662 2466 14714
rect 2466 14662 2478 14714
rect 2478 14662 2492 14714
rect 2516 14662 2530 14714
rect 2530 14662 2542 14714
rect 2542 14662 2572 14714
rect 2596 14662 2606 14714
rect 2606 14662 2652 14714
rect 2356 14660 2412 14662
rect 2436 14660 2492 14662
rect 2516 14660 2572 14662
rect 2596 14660 2652 14662
rect 3016 14170 3072 14172
rect 3096 14170 3152 14172
rect 3176 14170 3232 14172
rect 3256 14170 3312 14172
rect 3016 14118 3062 14170
rect 3062 14118 3072 14170
rect 3096 14118 3126 14170
rect 3126 14118 3138 14170
rect 3138 14118 3152 14170
rect 3176 14118 3190 14170
rect 3190 14118 3202 14170
rect 3202 14118 3232 14170
rect 3256 14118 3266 14170
rect 3266 14118 3312 14170
rect 3016 14116 3072 14118
rect 3096 14116 3152 14118
rect 3176 14116 3232 14118
rect 3256 14116 3312 14118
rect 2356 13626 2412 13628
rect 2436 13626 2492 13628
rect 2516 13626 2572 13628
rect 2596 13626 2652 13628
rect 2356 13574 2402 13626
rect 2402 13574 2412 13626
rect 2436 13574 2466 13626
rect 2466 13574 2478 13626
rect 2478 13574 2492 13626
rect 2516 13574 2530 13626
rect 2530 13574 2542 13626
rect 2542 13574 2572 13626
rect 2596 13574 2606 13626
rect 2606 13574 2652 13626
rect 2356 13572 2412 13574
rect 2436 13572 2492 13574
rect 2516 13572 2572 13574
rect 2596 13572 2652 13574
rect 1674 12280 1730 12336
rect 3016 13082 3072 13084
rect 3096 13082 3152 13084
rect 3176 13082 3232 13084
rect 3256 13082 3312 13084
rect 3016 13030 3062 13082
rect 3062 13030 3072 13082
rect 3096 13030 3126 13082
rect 3126 13030 3138 13082
rect 3138 13030 3152 13082
rect 3176 13030 3190 13082
rect 3190 13030 3202 13082
rect 3202 13030 3232 13082
rect 3256 13030 3266 13082
rect 3266 13030 3312 13082
rect 3016 13028 3072 13030
rect 3096 13028 3152 13030
rect 3176 13028 3232 13030
rect 3256 13028 3312 13030
rect 2356 12538 2412 12540
rect 2436 12538 2492 12540
rect 2516 12538 2572 12540
rect 2596 12538 2652 12540
rect 2356 12486 2402 12538
rect 2402 12486 2412 12538
rect 2436 12486 2466 12538
rect 2466 12486 2478 12538
rect 2478 12486 2492 12538
rect 2516 12486 2530 12538
rect 2530 12486 2542 12538
rect 2542 12486 2572 12538
rect 2596 12486 2606 12538
rect 2606 12486 2652 12538
rect 2356 12484 2412 12486
rect 2436 12484 2492 12486
rect 2516 12484 2572 12486
rect 2596 12484 2652 12486
rect 3016 11994 3072 11996
rect 3096 11994 3152 11996
rect 3176 11994 3232 11996
rect 3256 11994 3312 11996
rect 3016 11942 3062 11994
rect 3062 11942 3072 11994
rect 3096 11942 3126 11994
rect 3126 11942 3138 11994
rect 3138 11942 3152 11994
rect 3176 11942 3190 11994
rect 3190 11942 3202 11994
rect 3202 11942 3232 11994
rect 3256 11942 3266 11994
rect 3266 11942 3312 11994
rect 3016 11940 3072 11942
rect 3096 11940 3152 11942
rect 3176 11940 3232 11942
rect 3256 11940 3312 11942
rect 2356 11450 2412 11452
rect 2436 11450 2492 11452
rect 2516 11450 2572 11452
rect 2596 11450 2652 11452
rect 2356 11398 2402 11450
rect 2402 11398 2412 11450
rect 2436 11398 2466 11450
rect 2466 11398 2478 11450
rect 2478 11398 2492 11450
rect 2516 11398 2530 11450
rect 2530 11398 2542 11450
rect 2542 11398 2572 11450
rect 2596 11398 2606 11450
rect 2606 11398 2652 11450
rect 2356 11396 2412 11398
rect 2436 11396 2492 11398
rect 2516 11396 2572 11398
rect 2596 11396 2652 11398
rect 1398 10920 1454 10976
rect 17498 21800 17554 21856
rect 3790 11600 3846 11656
rect 846 10124 902 10160
rect 846 10104 848 10124
rect 848 10104 900 10124
rect 900 10104 902 10124
rect 2356 10362 2412 10364
rect 2436 10362 2492 10364
rect 2516 10362 2572 10364
rect 2596 10362 2652 10364
rect 2356 10310 2402 10362
rect 2402 10310 2412 10362
rect 2436 10310 2466 10362
rect 2466 10310 2478 10362
rect 2478 10310 2492 10362
rect 2516 10310 2530 10362
rect 2530 10310 2542 10362
rect 2542 10310 2572 10362
rect 2596 10310 2606 10362
rect 2606 10310 2652 10362
rect 2356 10308 2412 10310
rect 2436 10308 2492 10310
rect 2516 10308 2572 10310
rect 2596 10308 2652 10310
rect 846 9424 902 9480
rect 846 9052 848 9072
rect 848 9052 900 9072
rect 900 9052 902 9072
rect 846 9016 902 9052
rect 2356 9274 2412 9276
rect 2436 9274 2492 9276
rect 2516 9274 2572 9276
rect 2596 9274 2652 9276
rect 2356 9222 2402 9274
rect 2402 9222 2412 9274
rect 2436 9222 2466 9274
rect 2466 9222 2478 9274
rect 2478 9222 2492 9274
rect 2516 9222 2530 9274
rect 2530 9222 2542 9274
rect 2542 9222 2572 9274
rect 2596 9222 2606 9274
rect 2606 9222 2652 9274
rect 2356 9220 2412 9222
rect 2436 9220 2492 9222
rect 2516 9220 2572 9222
rect 2596 9220 2652 9222
rect 1306 8200 1362 8256
rect 2356 8186 2412 8188
rect 2436 8186 2492 8188
rect 2516 8186 2572 8188
rect 2596 8186 2652 8188
rect 2356 8134 2402 8186
rect 2402 8134 2412 8186
rect 2436 8134 2466 8186
rect 2466 8134 2478 8186
rect 2478 8134 2492 8186
rect 2516 8134 2530 8186
rect 2530 8134 2542 8186
rect 2542 8134 2572 8186
rect 2596 8134 2606 8186
rect 2606 8134 2652 8186
rect 2356 8132 2412 8134
rect 2436 8132 2492 8134
rect 2516 8132 2572 8134
rect 2596 8132 2652 8134
rect 1306 7540 1362 7576
rect 1306 7520 1308 7540
rect 1308 7520 1360 7540
rect 1360 7520 1362 7540
rect 2356 7098 2412 7100
rect 2436 7098 2492 7100
rect 2516 7098 2572 7100
rect 2596 7098 2652 7100
rect 2356 7046 2402 7098
rect 2402 7046 2412 7098
rect 2436 7046 2466 7098
rect 2466 7046 2478 7098
rect 2478 7046 2492 7098
rect 2516 7046 2530 7098
rect 2530 7046 2542 7098
rect 2542 7046 2572 7098
rect 2596 7046 2606 7098
rect 2606 7046 2652 7098
rect 2356 7044 2412 7046
rect 2436 7044 2492 7046
rect 2516 7044 2572 7046
rect 2596 7044 2652 7046
rect 846 6024 902 6080
rect 1490 5516 1492 5536
rect 1492 5516 1544 5536
rect 1544 5516 1546 5536
rect 1490 5480 1546 5516
rect 3016 10906 3072 10908
rect 3096 10906 3152 10908
rect 3176 10906 3232 10908
rect 3256 10906 3312 10908
rect 3016 10854 3062 10906
rect 3062 10854 3072 10906
rect 3096 10854 3126 10906
rect 3126 10854 3138 10906
rect 3138 10854 3152 10906
rect 3176 10854 3190 10906
rect 3190 10854 3202 10906
rect 3202 10854 3232 10906
rect 3256 10854 3266 10906
rect 3266 10854 3312 10906
rect 3016 10852 3072 10854
rect 3096 10852 3152 10854
rect 3176 10852 3232 10854
rect 3256 10852 3312 10854
rect 3016 9818 3072 9820
rect 3096 9818 3152 9820
rect 3176 9818 3232 9820
rect 3256 9818 3312 9820
rect 3016 9766 3062 9818
rect 3062 9766 3072 9818
rect 3096 9766 3126 9818
rect 3126 9766 3138 9818
rect 3138 9766 3152 9818
rect 3176 9766 3190 9818
rect 3190 9766 3202 9818
rect 3202 9766 3232 9818
rect 3256 9766 3266 9818
rect 3266 9766 3312 9818
rect 3016 9764 3072 9766
rect 3096 9764 3152 9766
rect 3176 9764 3232 9766
rect 3256 9764 3312 9766
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 1582 4800 1638 4856
rect 846 4256 902 4312
rect 846 3576 902 3632
rect 2356 6010 2412 6012
rect 2436 6010 2492 6012
rect 2516 6010 2572 6012
rect 2596 6010 2652 6012
rect 2356 5958 2402 6010
rect 2402 5958 2412 6010
rect 2436 5958 2466 6010
rect 2466 5958 2478 6010
rect 2478 5958 2492 6010
rect 2516 5958 2530 6010
rect 2530 5958 2542 6010
rect 2542 5958 2572 6010
rect 2596 5958 2606 6010
rect 2606 5958 2652 6010
rect 2356 5956 2412 5958
rect 2436 5956 2492 5958
rect 2516 5956 2572 5958
rect 2596 5956 2652 5958
rect 2356 4922 2412 4924
rect 2436 4922 2492 4924
rect 2516 4922 2572 4924
rect 2596 4922 2652 4924
rect 2356 4870 2402 4922
rect 2402 4870 2412 4922
rect 2436 4870 2466 4922
rect 2466 4870 2478 4922
rect 2478 4870 2492 4922
rect 2516 4870 2530 4922
rect 2530 4870 2542 4922
rect 2542 4870 2572 4922
rect 2596 4870 2606 4922
rect 2606 4870 2652 4922
rect 2356 4868 2412 4870
rect 2436 4868 2492 4870
rect 2516 4868 2572 4870
rect 2596 4868 2652 4870
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 17774 21120 17830 21176
rect 17958 20440 18014 20496
rect 16578 17720 16634 17776
rect 17590 17040 17646 17096
rect 4066 6704 4122 6760
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 2356 3834 2412 3836
rect 2436 3834 2492 3836
rect 2516 3834 2572 3836
rect 2596 3834 2652 3836
rect 2356 3782 2402 3834
rect 2402 3782 2412 3834
rect 2436 3782 2466 3834
rect 2466 3782 2478 3834
rect 2478 3782 2492 3834
rect 2516 3782 2530 3834
rect 2530 3782 2542 3834
rect 2542 3782 2572 3834
rect 2596 3782 2606 3834
rect 2606 3782 2652 3834
rect 2356 3780 2412 3782
rect 2436 3780 2492 3782
rect 2516 3780 2572 3782
rect 2596 3780 2652 3782
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 846 2896 902 2952
rect 2356 2746 2412 2748
rect 2436 2746 2492 2748
rect 2516 2746 2572 2748
rect 2596 2746 2652 2748
rect 2356 2694 2402 2746
rect 2402 2694 2412 2746
rect 2436 2694 2466 2746
rect 2466 2694 2478 2746
rect 2478 2694 2492 2746
rect 2516 2694 2530 2746
rect 2530 2694 2542 2746
rect 2542 2694 2572 2746
rect 2596 2694 2606 2746
rect 2606 2694 2652 2746
rect 2356 2692 2412 2694
rect 2436 2692 2492 2694
rect 2516 2692 2572 2694
rect 2596 2692 2652 2694
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 17498 11600 17554 11656
rect 18050 19760 18106 19816
rect 18050 19080 18106 19136
rect 18786 18420 18842 18456
rect 18786 18400 18788 18420
rect 18788 18400 18840 18420
rect 18840 18400 18842 18420
rect 18786 16360 18842 16416
rect 18786 15680 18842 15736
rect 18786 15000 18842 15056
rect 18878 14320 18934 14376
rect 18786 13640 18842 13696
rect 18786 12960 18842 13016
rect 18786 12280 18842 12336
rect 17406 8200 17462 8256
rect 18786 10920 18842 10976
rect 18786 10240 18842 10296
rect 18786 9560 18842 9616
rect 18510 8880 18566 8936
rect 17590 4800 17646 4856
rect 18786 7520 18842 7576
rect 18786 6840 18842 6896
rect 18786 6160 18842 6216
rect 18786 5480 18842 5536
rect 17682 1400 17738 1456
rect 18786 4120 18842 4176
rect 18786 3440 18842 3496
rect 18510 2760 18566 2816
rect 18142 2080 18198 2136
rect 17958 720 18014 776
rect 18234 40 18290 96
<< metal3 >>
rect 17493 21858 17559 21861
rect 19457 21858 20257 21888
rect 17493 21856 20257 21858
rect 17493 21800 17498 21856
rect 17554 21800 20257 21856
rect 17493 21798 20257 21800
rect 17493 21795 17559 21798
rect 19457 21768 20257 21798
rect 17769 21178 17835 21181
rect 19457 21178 20257 21208
rect 17769 21176 20257 21178
rect 17769 21120 17774 21176
rect 17830 21120 20257 21176
rect 17769 21118 20257 21120
rect 17769 21115 17835 21118
rect 19457 21088 20257 21118
rect 17953 20498 18019 20501
rect 19457 20498 20257 20528
rect 17953 20496 20257 20498
rect 17953 20440 17958 20496
rect 18014 20440 20257 20496
rect 17953 20438 20257 20440
rect 17953 20435 18019 20438
rect 19457 20408 20257 20438
rect 2346 20160 2662 20161
rect 2346 20096 2352 20160
rect 2416 20096 2432 20160
rect 2496 20096 2512 20160
rect 2576 20096 2592 20160
rect 2656 20096 2662 20160
rect 2346 20095 2662 20096
rect 18045 19818 18111 19821
rect 19457 19818 20257 19848
rect 18045 19816 20257 19818
rect 18045 19760 18050 19816
rect 18106 19760 20257 19816
rect 18045 19758 20257 19760
rect 18045 19755 18111 19758
rect 19457 19728 20257 19758
rect 3006 19616 3322 19617
rect 3006 19552 3012 19616
rect 3076 19552 3092 19616
rect 3156 19552 3172 19616
rect 3236 19552 3252 19616
rect 3316 19552 3322 19616
rect 3006 19551 3322 19552
rect 5073 19274 5139 19277
rect 2086 19272 5139 19274
rect 2086 19216 5078 19272
rect 5134 19216 5139 19272
rect 2086 19214 5139 19216
rect 0 19138 800 19168
rect 2086 19138 2146 19214
rect 5073 19211 5139 19214
rect 0 19078 2146 19138
rect 18045 19138 18111 19141
rect 19457 19138 20257 19168
rect 18045 19136 20257 19138
rect 18045 19080 18050 19136
rect 18106 19080 20257 19136
rect 18045 19078 20257 19080
rect 0 19048 800 19078
rect 18045 19075 18111 19078
rect 2346 19072 2662 19073
rect 2346 19008 2352 19072
rect 2416 19008 2432 19072
rect 2496 19008 2512 19072
rect 2576 19008 2592 19072
rect 2656 19008 2662 19072
rect 19457 19048 20257 19078
rect 2346 19007 2662 19008
rect 841 18594 907 18597
rect 798 18592 907 18594
rect 798 18536 846 18592
rect 902 18536 907 18592
rect 798 18531 907 18536
rect 798 18488 858 18531
rect 0 18398 858 18488
rect 3006 18528 3322 18529
rect 3006 18464 3012 18528
rect 3076 18464 3092 18528
rect 3156 18464 3172 18528
rect 3236 18464 3252 18528
rect 3316 18464 3322 18528
rect 3006 18463 3322 18464
rect 18781 18458 18847 18461
rect 19457 18458 20257 18488
rect 18781 18456 20257 18458
rect 18781 18400 18786 18456
rect 18842 18400 20257 18456
rect 18781 18398 20257 18400
rect 0 18368 800 18398
rect 18781 18395 18847 18398
rect 19457 18368 20257 18398
rect 2346 17984 2662 17985
rect 2346 17920 2352 17984
rect 2416 17920 2432 17984
rect 2496 17920 2512 17984
rect 2576 17920 2592 17984
rect 2656 17920 2662 17984
rect 2346 17919 2662 17920
rect 0 17778 800 17808
rect 16573 17778 16639 17781
rect 19457 17778 20257 17808
rect 0 17688 858 17778
rect 16573 17776 20257 17778
rect 16573 17720 16578 17776
rect 16634 17720 20257 17776
rect 16573 17718 20257 17720
rect 16573 17715 16639 17718
rect 19457 17688 20257 17718
rect 798 17645 858 17688
rect 798 17640 907 17645
rect 798 17584 846 17640
rect 902 17584 907 17640
rect 798 17582 907 17584
rect 841 17579 907 17582
rect 3006 17440 3322 17441
rect 3006 17376 3012 17440
rect 3076 17376 3092 17440
rect 3156 17376 3172 17440
rect 3236 17376 3252 17440
rect 3316 17376 3322 17440
rect 3006 17375 3322 17376
rect 0 17098 800 17128
rect 1209 17098 1275 17101
rect 0 17096 1275 17098
rect 0 17040 1214 17096
rect 1270 17040 1275 17096
rect 0 17038 1275 17040
rect 0 17008 800 17038
rect 1209 17035 1275 17038
rect 17585 17098 17651 17101
rect 19457 17098 20257 17128
rect 17585 17096 20257 17098
rect 17585 17040 17590 17096
rect 17646 17040 20257 17096
rect 17585 17038 20257 17040
rect 17585 17035 17651 17038
rect 19457 17008 20257 17038
rect 2346 16896 2662 16897
rect 2346 16832 2352 16896
rect 2416 16832 2432 16896
rect 2496 16832 2512 16896
rect 2576 16832 2592 16896
rect 2656 16832 2662 16896
rect 2346 16831 2662 16832
rect 0 16418 800 16448
rect 1393 16418 1459 16421
rect 0 16416 1459 16418
rect 0 16360 1398 16416
rect 1454 16360 1459 16416
rect 0 16358 1459 16360
rect 0 16328 800 16358
rect 1393 16355 1459 16358
rect 18781 16418 18847 16421
rect 19457 16418 20257 16448
rect 18781 16416 20257 16418
rect 18781 16360 18786 16416
rect 18842 16360 20257 16416
rect 18781 16358 20257 16360
rect 18781 16355 18847 16358
rect 3006 16352 3322 16353
rect 3006 16288 3012 16352
rect 3076 16288 3092 16352
rect 3156 16288 3172 16352
rect 3236 16288 3252 16352
rect 3316 16288 3322 16352
rect 19457 16328 20257 16358
rect 3006 16287 3322 16288
rect 841 15874 907 15877
rect 798 15872 907 15874
rect 798 15816 846 15872
rect 902 15816 907 15872
rect 798 15811 907 15816
rect 798 15768 858 15811
rect 0 15678 858 15768
rect 2346 15808 2662 15809
rect 2346 15744 2352 15808
rect 2416 15744 2432 15808
rect 2496 15744 2512 15808
rect 2576 15744 2592 15808
rect 2656 15744 2662 15808
rect 2346 15743 2662 15744
rect 18781 15738 18847 15741
rect 19457 15738 20257 15768
rect 18781 15736 20257 15738
rect 18781 15680 18786 15736
rect 18842 15680 20257 15736
rect 18781 15678 20257 15680
rect 0 15648 800 15678
rect 18781 15675 18847 15678
rect 19457 15648 20257 15678
rect 3006 15264 3322 15265
rect 3006 15200 3012 15264
rect 3076 15200 3092 15264
rect 3156 15200 3172 15264
rect 3236 15200 3252 15264
rect 3316 15200 3322 15264
rect 3006 15199 3322 15200
rect 0 15058 800 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 800 14998
rect 1393 14995 1459 14998
rect 18781 15058 18847 15061
rect 19457 15058 20257 15088
rect 18781 15056 20257 15058
rect 18781 15000 18786 15056
rect 18842 15000 20257 15056
rect 18781 14998 20257 15000
rect 18781 14995 18847 14998
rect 19457 14968 20257 14998
rect 2346 14720 2662 14721
rect 2346 14656 2352 14720
rect 2416 14656 2432 14720
rect 2496 14656 2512 14720
rect 2576 14656 2592 14720
rect 2656 14656 2662 14720
rect 2346 14655 2662 14656
rect 0 14378 800 14408
rect 1025 14378 1091 14381
rect 0 14376 1091 14378
rect 0 14320 1030 14376
rect 1086 14320 1091 14376
rect 0 14318 1091 14320
rect 0 14288 800 14318
rect 1025 14315 1091 14318
rect 18873 14378 18939 14381
rect 19457 14378 20257 14408
rect 18873 14376 20257 14378
rect 18873 14320 18878 14376
rect 18934 14320 20257 14376
rect 18873 14318 20257 14320
rect 18873 14315 18939 14318
rect 19457 14288 20257 14318
rect 3006 14176 3322 14177
rect 3006 14112 3012 14176
rect 3076 14112 3092 14176
rect 3156 14112 3172 14176
rect 3236 14112 3252 14176
rect 3316 14112 3322 14176
rect 3006 14111 3322 14112
rect 0 13698 800 13728
rect 1485 13698 1551 13701
rect 0 13696 1551 13698
rect 0 13640 1490 13696
rect 1546 13640 1551 13696
rect 0 13638 1551 13640
rect 0 13608 800 13638
rect 1485 13635 1551 13638
rect 18781 13698 18847 13701
rect 19457 13698 20257 13728
rect 18781 13696 20257 13698
rect 18781 13640 18786 13696
rect 18842 13640 20257 13696
rect 18781 13638 20257 13640
rect 18781 13635 18847 13638
rect 2346 13632 2662 13633
rect 2346 13568 2352 13632
rect 2416 13568 2432 13632
rect 2496 13568 2512 13632
rect 2576 13568 2592 13632
rect 2656 13568 2662 13632
rect 19457 13608 20257 13638
rect 2346 13567 2662 13568
rect 3006 13088 3322 13089
rect 0 13018 800 13048
rect 3006 13024 3012 13088
rect 3076 13024 3092 13088
rect 3156 13024 3172 13088
rect 3236 13024 3252 13088
rect 3316 13024 3322 13088
rect 3006 13023 3322 13024
rect 1209 13018 1275 13021
rect 0 13016 1275 13018
rect 0 12960 1214 13016
rect 1270 12960 1275 13016
rect 0 12958 1275 12960
rect 0 12928 800 12958
rect 1209 12955 1275 12958
rect 18781 13018 18847 13021
rect 19457 13018 20257 13048
rect 18781 13016 20257 13018
rect 18781 12960 18786 13016
rect 18842 12960 20257 13016
rect 18781 12958 20257 12960
rect 18781 12955 18847 12958
rect 19457 12928 20257 12958
rect 2346 12544 2662 12545
rect 2346 12480 2352 12544
rect 2416 12480 2432 12544
rect 2496 12480 2512 12544
rect 2576 12480 2592 12544
rect 2656 12480 2662 12544
rect 2346 12479 2662 12480
rect 0 12338 800 12368
rect 1669 12338 1735 12341
rect 0 12336 1735 12338
rect 0 12280 1674 12336
rect 1730 12280 1735 12336
rect 0 12278 1735 12280
rect 0 12248 800 12278
rect 1669 12275 1735 12278
rect 18781 12338 18847 12341
rect 19457 12338 20257 12368
rect 18781 12336 20257 12338
rect 18781 12280 18786 12336
rect 18842 12280 20257 12336
rect 18781 12278 20257 12280
rect 18781 12275 18847 12278
rect 19457 12248 20257 12278
rect 3006 12000 3322 12001
rect 3006 11936 3012 12000
rect 3076 11936 3092 12000
rect 3156 11936 3172 12000
rect 3236 11936 3252 12000
rect 3316 11936 3322 12000
rect 3006 11935 3322 11936
rect 0 11658 800 11688
rect 3785 11658 3851 11661
rect 0 11656 3851 11658
rect 0 11600 3790 11656
rect 3846 11600 3851 11656
rect 0 11598 3851 11600
rect 0 11568 800 11598
rect 3785 11595 3851 11598
rect 17493 11658 17559 11661
rect 19457 11658 20257 11688
rect 17493 11656 20257 11658
rect 17493 11600 17498 11656
rect 17554 11600 20257 11656
rect 17493 11598 20257 11600
rect 17493 11595 17559 11598
rect 19457 11568 20257 11598
rect 2346 11456 2662 11457
rect 2346 11392 2352 11456
rect 2416 11392 2432 11456
rect 2496 11392 2512 11456
rect 2576 11392 2592 11456
rect 2656 11392 2662 11456
rect 2346 11391 2662 11392
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 18781 10978 18847 10981
rect 19457 10978 20257 11008
rect 18781 10976 20257 10978
rect 18781 10920 18786 10976
rect 18842 10920 20257 10976
rect 18781 10918 20257 10920
rect 18781 10915 18847 10918
rect 3006 10912 3322 10913
rect 3006 10848 3012 10912
rect 3076 10848 3092 10912
rect 3156 10848 3172 10912
rect 3236 10848 3252 10912
rect 3316 10848 3322 10912
rect 19457 10888 20257 10918
rect 3006 10847 3322 10848
rect 2346 10368 2662 10369
rect 0 10298 800 10328
rect 2346 10304 2352 10368
rect 2416 10304 2432 10368
rect 2496 10304 2512 10368
rect 2576 10304 2592 10368
rect 2656 10304 2662 10368
rect 2346 10303 2662 10304
rect 18781 10298 18847 10301
rect 19457 10298 20257 10328
rect 0 10208 858 10298
rect 18781 10296 20257 10298
rect 18781 10240 18786 10296
rect 18842 10240 20257 10296
rect 18781 10238 20257 10240
rect 18781 10235 18847 10238
rect 19457 10208 20257 10238
rect 798 10165 858 10208
rect 798 10160 907 10165
rect 798 10104 846 10160
rect 902 10104 907 10160
rect 798 10102 907 10104
rect 841 10099 907 10102
rect 3006 9824 3322 9825
rect 3006 9760 3012 9824
rect 3076 9760 3092 9824
rect 3156 9760 3172 9824
rect 3236 9760 3252 9824
rect 3316 9760 3322 9824
rect 3006 9759 3322 9760
rect 0 9618 800 9648
rect 18781 9618 18847 9621
rect 19457 9618 20257 9648
rect 0 9528 858 9618
rect 18781 9616 20257 9618
rect 18781 9560 18786 9616
rect 18842 9560 20257 9616
rect 18781 9558 20257 9560
rect 18781 9555 18847 9558
rect 19457 9528 20257 9558
rect 798 9485 858 9528
rect 798 9480 907 9485
rect 798 9424 846 9480
rect 902 9424 907 9480
rect 798 9422 907 9424
rect 841 9419 907 9422
rect 2346 9280 2662 9281
rect 2346 9216 2352 9280
rect 2416 9216 2432 9280
rect 2496 9216 2512 9280
rect 2576 9216 2592 9280
rect 2656 9216 2662 9280
rect 2346 9215 2662 9216
rect 841 9074 907 9077
rect 798 9072 907 9074
rect 798 9016 846 9072
rect 902 9016 907 9072
rect 798 9011 907 9016
rect 798 8968 858 9011
rect 0 8878 858 8968
rect 18505 8938 18571 8941
rect 19457 8938 20257 8968
rect 18505 8936 20257 8938
rect 18505 8880 18510 8936
rect 18566 8880 20257 8936
rect 18505 8878 20257 8880
rect 0 8848 800 8878
rect 18505 8875 18571 8878
rect 19457 8848 20257 8878
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 0 8258 800 8288
rect 1301 8258 1367 8261
rect 0 8256 1367 8258
rect 0 8200 1306 8256
rect 1362 8200 1367 8256
rect 0 8198 1367 8200
rect 0 8168 800 8198
rect 1301 8195 1367 8198
rect 17401 8258 17467 8261
rect 19457 8258 20257 8288
rect 17401 8256 20257 8258
rect 17401 8200 17406 8256
rect 17462 8200 20257 8256
rect 17401 8198 20257 8200
rect 17401 8195 17467 8198
rect 2346 8192 2662 8193
rect 2346 8128 2352 8192
rect 2416 8128 2432 8192
rect 2496 8128 2512 8192
rect 2576 8128 2592 8192
rect 2656 8128 2662 8192
rect 19457 8168 20257 8198
rect 2346 8127 2662 8128
rect 3006 7648 3322 7649
rect 0 7578 800 7608
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 1301 7578 1367 7581
rect 0 7576 1367 7578
rect 0 7520 1306 7576
rect 1362 7520 1367 7576
rect 0 7518 1367 7520
rect 0 7488 800 7518
rect 1301 7515 1367 7518
rect 18781 7578 18847 7581
rect 19457 7578 20257 7608
rect 18781 7576 20257 7578
rect 18781 7520 18786 7576
rect 18842 7520 20257 7576
rect 18781 7518 20257 7520
rect 18781 7515 18847 7518
rect 19457 7488 20257 7518
rect 2346 7104 2662 7105
rect 2346 7040 2352 7104
rect 2416 7040 2432 7104
rect 2496 7040 2512 7104
rect 2576 7040 2592 7104
rect 2656 7040 2662 7104
rect 2346 7039 2662 7040
rect 0 6898 800 6928
rect 18781 6898 18847 6901
rect 19457 6898 20257 6928
rect 0 6838 2790 6898
rect 0 6808 800 6838
rect 2730 6762 2790 6838
rect 18781 6896 20257 6898
rect 18781 6840 18786 6896
rect 18842 6840 20257 6896
rect 18781 6838 20257 6840
rect 18781 6835 18847 6838
rect 19457 6808 20257 6838
rect 4061 6762 4127 6765
rect 2730 6760 4127 6762
rect 2730 6704 4066 6760
rect 4122 6704 4127 6760
rect 2730 6702 4127 6704
rect 4061 6699 4127 6702
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 0 6218 800 6248
rect 18781 6218 18847 6221
rect 19457 6218 20257 6248
rect 0 6128 858 6218
rect 18781 6216 20257 6218
rect 18781 6160 18786 6216
rect 18842 6160 20257 6216
rect 18781 6158 20257 6160
rect 18781 6155 18847 6158
rect 19457 6128 20257 6158
rect 798 6085 858 6128
rect 798 6080 907 6085
rect 798 6024 846 6080
rect 902 6024 907 6080
rect 798 6022 907 6024
rect 841 6019 907 6022
rect 2346 6016 2662 6017
rect 2346 5952 2352 6016
rect 2416 5952 2432 6016
rect 2496 5952 2512 6016
rect 2576 5952 2592 6016
rect 2656 5952 2662 6016
rect 2346 5951 2662 5952
rect 0 5538 800 5568
rect 1485 5538 1551 5541
rect 0 5536 1551 5538
rect 0 5480 1490 5536
rect 1546 5480 1551 5536
rect 0 5478 1551 5480
rect 0 5448 800 5478
rect 1485 5475 1551 5478
rect 18781 5538 18847 5541
rect 19457 5538 20257 5568
rect 18781 5536 20257 5538
rect 18781 5480 18786 5536
rect 18842 5480 20257 5536
rect 18781 5478 20257 5480
rect 18781 5475 18847 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 19457 5448 20257 5478
rect 3006 5407 3322 5408
rect 2346 4928 2662 4929
rect 0 4858 800 4888
rect 2346 4864 2352 4928
rect 2416 4864 2432 4928
rect 2496 4864 2512 4928
rect 2576 4864 2592 4928
rect 2656 4864 2662 4928
rect 2346 4863 2662 4864
rect 1577 4858 1643 4861
rect 0 4856 1643 4858
rect 0 4800 1582 4856
rect 1638 4800 1643 4856
rect 0 4798 1643 4800
rect 0 4768 800 4798
rect 1577 4795 1643 4798
rect 17585 4858 17651 4861
rect 19457 4858 20257 4888
rect 17585 4856 20257 4858
rect 17585 4800 17590 4856
rect 17646 4800 20257 4856
rect 17585 4798 20257 4800
rect 17585 4795 17651 4798
rect 19457 4768 20257 4798
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 841 4314 907 4317
rect 798 4312 907 4314
rect 798 4256 846 4312
rect 902 4256 907 4312
rect 798 4251 907 4256
rect 798 4208 858 4251
rect 0 4118 858 4208
rect 18781 4178 18847 4181
rect 19457 4178 20257 4208
rect 18781 4176 20257 4178
rect 18781 4120 18786 4176
rect 18842 4120 20257 4176
rect 18781 4118 20257 4120
rect 0 4088 800 4118
rect 18781 4115 18847 4118
rect 19457 4088 20257 4118
rect 2346 3840 2662 3841
rect 2346 3776 2352 3840
rect 2416 3776 2432 3840
rect 2496 3776 2512 3840
rect 2576 3776 2592 3840
rect 2656 3776 2662 3840
rect 2346 3775 2662 3776
rect 841 3634 907 3637
rect 798 3632 907 3634
rect 798 3576 846 3632
rect 902 3576 907 3632
rect 798 3571 907 3576
rect 798 3528 858 3571
rect 0 3438 858 3528
rect 18781 3498 18847 3501
rect 19457 3498 20257 3528
rect 18781 3496 20257 3498
rect 18781 3440 18786 3496
rect 18842 3440 20257 3496
rect 18781 3438 20257 3440
rect 0 3408 800 3438
rect 18781 3435 18847 3438
rect 19457 3408 20257 3438
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 841 2954 907 2957
rect 798 2952 907 2954
rect 798 2896 846 2952
rect 902 2896 907 2952
rect 798 2891 907 2896
rect 798 2848 858 2891
rect 0 2758 858 2848
rect 18505 2818 18571 2821
rect 19457 2818 20257 2848
rect 18505 2816 20257 2818
rect 18505 2760 18510 2816
rect 18566 2760 20257 2816
rect 18505 2758 20257 2760
rect 0 2728 800 2758
rect 18505 2755 18571 2758
rect 2346 2752 2662 2753
rect 2346 2688 2352 2752
rect 2416 2688 2432 2752
rect 2496 2688 2512 2752
rect 2576 2688 2592 2752
rect 2656 2688 2662 2752
rect 19457 2728 20257 2758
rect 2346 2687 2662 2688
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 18137 2138 18203 2141
rect 19457 2138 20257 2168
rect 18137 2136 20257 2138
rect 18137 2080 18142 2136
rect 18198 2080 20257 2136
rect 18137 2078 20257 2080
rect 18137 2075 18203 2078
rect 19457 2048 20257 2078
rect 17677 1458 17743 1461
rect 19457 1458 20257 1488
rect 17677 1456 20257 1458
rect 17677 1400 17682 1456
rect 17738 1400 20257 1456
rect 17677 1398 20257 1400
rect 17677 1395 17743 1398
rect 19457 1368 20257 1398
rect 17953 778 18019 781
rect 19457 778 20257 808
rect 17953 776 20257 778
rect 17953 720 17958 776
rect 18014 720 20257 776
rect 17953 718 20257 720
rect 17953 715 18019 718
rect 19457 688 20257 718
rect 18229 98 18295 101
rect 19457 98 20257 128
rect 18229 96 20257 98
rect 18229 40 18234 96
rect 18290 40 20257 96
rect 18229 38 20257 40
rect 18229 35 18295 38
rect 19457 8 20257 38
<< via3 >>
rect 2352 20156 2416 20160
rect 2352 20100 2356 20156
rect 2356 20100 2412 20156
rect 2412 20100 2416 20156
rect 2352 20096 2416 20100
rect 2432 20156 2496 20160
rect 2432 20100 2436 20156
rect 2436 20100 2492 20156
rect 2492 20100 2496 20156
rect 2432 20096 2496 20100
rect 2512 20156 2576 20160
rect 2512 20100 2516 20156
rect 2516 20100 2572 20156
rect 2572 20100 2576 20156
rect 2512 20096 2576 20100
rect 2592 20156 2656 20160
rect 2592 20100 2596 20156
rect 2596 20100 2652 20156
rect 2652 20100 2656 20156
rect 2592 20096 2656 20100
rect 3012 19612 3076 19616
rect 3012 19556 3016 19612
rect 3016 19556 3072 19612
rect 3072 19556 3076 19612
rect 3012 19552 3076 19556
rect 3092 19612 3156 19616
rect 3092 19556 3096 19612
rect 3096 19556 3152 19612
rect 3152 19556 3156 19612
rect 3092 19552 3156 19556
rect 3172 19612 3236 19616
rect 3172 19556 3176 19612
rect 3176 19556 3232 19612
rect 3232 19556 3236 19612
rect 3172 19552 3236 19556
rect 3252 19612 3316 19616
rect 3252 19556 3256 19612
rect 3256 19556 3312 19612
rect 3312 19556 3316 19612
rect 3252 19552 3316 19556
rect 2352 19068 2416 19072
rect 2352 19012 2356 19068
rect 2356 19012 2412 19068
rect 2412 19012 2416 19068
rect 2352 19008 2416 19012
rect 2432 19068 2496 19072
rect 2432 19012 2436 19068
rect 2436 19012 2492 19068
rect 2492 19012 2496 19068
rect 2432 19008 2496 19012
rect 2512 19068 2576 19072
rect 2512 19012 2516 19068
rect 2516 19012 2572 19068
rect 2572 19012 2576 19068
rect 2512 19008 2576 19012
rect 2592 19068 2656 19072
rect 2592 19012 2596 19068
rect 2596 19012 2652 19068
rect 2652 19012 2656 19068
rect 2592 19008 2656 19012
rect 3012 18524 3076 18528
rect 3012 18468 3016 18524
rect 3016 18468 3072 18524
rect 3072 18468 3076 18524
rect 3012 18464 3076 18468
rect 3092 18524 3156 18528
rect 3092 18468 3096 18524
rect 3096 18468 3152 18524
rect 3152 18468 3156 18524
rect 3092 18464 3156 18468
rect 3172 18524 3236 18528
rect 3172 18468 3176 18524
rect 3176 18468 3232 18524
rect 3232 18468 3236 18524
rect 3172 18464 3236 18468
rect 3252 18524 3316 18528
rect 3252 18468 3256 18524
rect 3256 18468 3312 18524
rect 3312 18468 3316 18524
rect 3252 18464 3316 18468
rect 2352 17980 2416 17984
rect 2352 17924 2356 17980
rect 2356 17924 2412 17980
rect 2412 17924 2416 17980
rect 2352 17920 2416 17924
rect 2432 17980 2496 17984
rect 2432 17924 2436 17980
rect 2436 17924 2492 17980
rect 2492 17924 2496 17980
rect 2432 17920 2496 17924
rect 2512 17980 2576 17984
rect 2512 17924 2516 17980
rect 2516 17924 2572 17980
rect 2572 17924 2576 17980
rect 2512 17920 2576 17924
rect 2592 17980 2656 17984
rect 2592 17924 2596 17980
rect 2596 17924 2652 17980
rect 2652 17924 2656 17980
rect 2592 17920 2656 17924
rect 3012 17436 3076 17440
rect 3012 17380 3016 17436
rect 3016 17380 3072 17436
rect 3072 17380 3076 17436
rect 3012 17376 3076 17380
rect 3092 17436 3156 17440
rect 3092 17380 3096 17436
rect 3096 17380 3152 17436
rect 3152 17380 3156 17436
rect 3092 17376 3156 17380
rect 3172 17436 3236 17440
rect 3172 17380 3176 17436
rect 3176 17380 3232 17436
rect 3232 17380 3236 17436
rect 3172 17376 3236 17380
rect 3252 17436 3316 17440
rect 3252 17380 3256 17436
rect 3256 17380 3312 17436
rect 3312 17380 3316 17436
rect 3252 17376 3316 17380
rect 2352 16892 2416 16896
rect 2352 16836 2356 16892
rect 2356 16836 2412 16892
rect 2412 16836 2416 16892
rect 2352 16832 2416 16836
rect 2432 16892 2496 16896
rect 2432 16836 2436 16892
rect 2436 16836 2492 16892
rect 2492 16836 2496 16892
rect 2432 16832 2496 16836
rect 2512 16892 2576 16896
rect 2512 16836 2516 16892
rect 2516 16836 2572 16892
rect 2572 16836 2576 16892
rect 2512 16832 2576 16836
rect 2592 16892 2656 16896
rect 2592 16836 2596 16892
rect 2596 16836 2652 16892
rect 2652 16836 2656 16892
rect 2592 16832 2656 16836
rect 3012 16348 3076 16352
rect 3012 16292 3016 16348
rect 3016 16292 3072 16348
rect 3072 16292 3076 16348
rect 3012 16288 3076 16292
rect 3092 16348 3156 16352
rect 3092 16292 3096 16348
rect 3096 16292 3152 16348
rect 3152 16292 3156 16348
rect 3092 16288 3156 16292
rect 3172 16348 3236 16352
rect 3172 16292 3176 16348
rect 3176 16292 3232 16348
rect 3232 16292 3236 16348
rect 3172 16288 3236 16292
rect 3252 16348 3316 16352
rect 3252 16292 3256 16348
rect 3256 16292 3312 16348
rect 3312 16292 3316 16348
rect 3252 16288 3316 16292
rect 2352 15804 2416 15808
rect 2352 15748 2356 15804
rect 2356 15748 2412 15804
rect 2412 15748 2416 15804
rect 2352 15744 2416 15748
rect 2432 15804 2496 15808
rect 2432 15748 2436 15804
rect 2436 15748 2492 15804
rect 2492 15748 2496 15804
rect 2432 15744 2496 15748
rect 2512 15804 2576 15808
rect 2512 15748 2516 15804
rect 2516 15748 2572 15804
rect 2572 15748 2576 15804
rect 2512 15744 2576 15748
rect 2592 15804 2656 15808
rect 2592 15748 2596 15804
rect 2596 15748 2652 15804
rect 2652 15748 2656 15804
rect 2592 15744 2656 15748
rect 3012 15260 3076 15264
rect 3012 15204 3016 15260
rect 3016 15204 3072 15260
rect 3072 15204 3076 15260
rect 3012 15200 3076 15204
rect 3092 15260 3156 15264
rect 3092 15204 3096 15260
rect 3096 15204 3152 15260
rect 3152 15204 3156 15260
rect 3092 15200 3156 15204
rect 3172 15260 3236 15264
rect 3172 15204 3176 15260
rect 3176 15204 3232 15260
rect 3232 15204 3236 15260
rect 3172 15200 3236 15204
rect 3252 15260 3316 15264
rect 3252 15204 3256 15260
rect 3256 15204 3312 15260
rect 3312 15204 3316 15260
rect 3252 15200 3316 15204
rect 2352 14716 2416 14720
rect 2352 14660 2356 14716
rect 2356 14660 2412 14716
rect 2412 14660 2416 14716
rect 2352 14656 2416 14660
rect 2432 14716 2496 14720
rect 2432 14660 2436 14716
rect 2436 14660 2492 14716
rect 2492 14660 2496 14716
rect 2432 14656 2496 14660
rect 2512 14716 2576 14720
rect 2512 14660 2516 14716
rect 2516 14660 2572 14716
rect 2572 14660 2576 14716
rect 2512 14656 2576 14660
rect 2592 14716 2656 14720
rect 2592 14660 2596 14716
rect 2596 14660 2652 14716
rect 2652 14660 2656 14716
rect 2592 14656 2656 14660
rect 3012 14172 3076 14176
rect 3012 14116 3016 14172
rect 3016 14116 3072 14172
rect 3072 14116 3076 14172
rect 3012 14112 3076 14116
rect 3092 14172 3156 14176
rect 3092 14116 3096 14172
rect 3096 14116 3152 14172
rect 3152 14116 3156 14172
rect 3092 14112 3156 14116
rect 3172 14172 3236 14176
rect 3172 14116 3176 14172
rect 3176 14116 3232 14172
rect 3232 14116 3236 14172
rect 3172 14112 3236 14116
rect 3252 14172 3316 14176
rect 3252 14116 3256 14172
rect 3256 14116 3312 14172
rect 3312 14116 3316 14172
rect 3252 14112 3316 14116
rect 2352 13628 2416 13632
rect 2352 13572 2356 13628
rect 2356 13572 2412 13628
rect 2412 13572 2416 13628
rect 2352 13568 2416 13572
rect 2432 13628 2496 13632
rect 2432 13572 2436 13628
rect 2436 13572 2492 13628
rect 2492 13572 2496 13628
rect 2432 13568 2496 13572
rect 2512 13628 2576 13632
rect 2512 13572 2516 13628
rect 2516 13572 2572 13628
rect 2572 13572 2576 13628
rect 2512 13568 2576 13572
rect 2592 13628 2656 13632
rect 2592 13572 2596 13628
rect 2596 13572 2652 13628
rect 2652 13572 2656 13628
rect 2592 13568 2656 13572
rect 3012 13084 3076 13088
rect 3012 13028 3016 13084
rect 3016 13028 3072 13084
rect 3072 13028 3076 13084
rect 3012 13024 3076 13028
rect 3092 13084 3156 13088
rect 3092 13028 3096 13084
rect 3096 13028 3152 13084
rect 3152 13028 3156 13084
rect 3092 13024 3156 13028
rect 3172 13084 3236 13088
rect 3172 13028 3176 13084
rect 3176 13028 3232 13084
rect 3232 13028 3236 13084
rect 3172 13024 3236 13028
rect 3252 13084 3316 13088
rect 3252 13028 3256 13084
rect 3256 13028 3312 13084
rect 3312 13028 3316 13084
rect 3252 13024 3316 13028
rect 2352 12540 2416 12544
rect 2352 12484 2356 12540
rect 2356 12484 2412 12540
rect 2412 12484 2416 12540
rect 2352 12480 2416 12484
rect 2432 12540 2496 12544
rect 2432 12484 2436 12540
rect 2436 12484 2492 12540
rect 2492 12484 2496 12540
rect 2432 12480 2496 12484
rect 2512 12540 2576 12544
rect 2512 12484 2516 12540
rect 2516 12484 2572 12540
rect 2572 12484 2576 12540
rect 2512 12480 2576 12484
rect 2592 12540 2656 12544
rect 2592 12484 2596 12540
rect 2596 12484 2652 12540
rect 2652 12484 2656 12540
rect 2592 12480 2656 12484
rect 3012 11996 3076 12000
rect 3012 11940 3016 11996
rect 3016 11940 3072 11996
rect 3072 11940 3076 11996
rect 3012 11936 3076 11940
rect 3092 11996 3156 12000
rect 3092 11940 3096 11996
rect 3096 11940 3152 11996
rect 3152 11940 3156 11996
rect 3092 11936 3156 11940
rect 3172 11996 3236 12000
rect 3172 11940 3176 11996
rect 3176 11940 3232 11996
rect 3232 11940 3236 11996
rect 3172 11936 3236 11940
rect 3252 11996 3316 12000
rect 3252 11940 3256 11996
rect 3256 11940 3312 11996
rect 3312 11940 3316 11996
rect 3252 11936 3316 11940
rect 2352 11452 2416 11456
rect 2352 11396 2356 11452
rect 2356 11396 2412 11452
rect 2412 11396 2416 11452
rect 2352 11392 2416 11396
rect 2432 11452 2496 11456
rect 2432 11396 2436 11452
rect 2436 11396 2492 11452
rect 2492 11396 2496 11452
rect 2432 11392 2496 11396
rect 2512 11452 2576 11456
rect 2512 11396 2516 11452
rect 2516 11396 2572 11452
rect 2572 11396 2576 11452
rect 2512 11392 2576 11396
rect 2592 11452 2656 11456
rect 2592 11396 2596 11452
rect 2596 11396 2652 11452
rect 2652 11396 2656 11452
rect 2592 11392 2656 11396
rect 3012 10908 3076 10912
rect 3012 10852 3016 10908
rect 3016 10852 3072 10908
rect 3072 10852 3076 10908
rect 3012 10848 3076 10852
rect 3092 10908 3156 10912
rect 3092 10852 3096 10908
rect 3096 10852 3152 10908
rect 3152 10852 3156 10908
rect 3092 10848 3156 10852
rect 3172 10908 3236 10912
rect 3172 10852 3176 10908
rect 3176 10852 3232 10908
rect 3232 10852 3236 10908
rect 3172 10848 3236 10852
rect 3252 10908 3316 10912
rect 3252 10852 3256 10908
rect 3256 10852 3312 10908
rect 3312 10852 3316 10908
rect 3252 10848 3316 10852
rect 2352 10364 2416 10368
rect 2352 10308 2356 10364
rect 2356 10308 2412 10364
rect 2412 10308 2416 10364
rect 2352 10304 2416 10308
rect 2432 10364 2496 10368
rect 2432 10308 2436 10364
rect 2436 10308 2492 10364
rect 2492 10308 2496 10364
rect 2432 10304 2496 10308
rect 2512 10364 2576 10368
rect 2512 10308 2516 10364
rect 2516 10308 2572 10364
rect 2572 10308 2576 10364
rect 2512 10304 2576 10308
rect 2592 10364 2656 10368
rect 2592 10308 2596 10364
rect 2596 10308 2652 10364
rect 2652 10308 2656 10364
rect 2592 10304 2656 10308
rect 3012 9820 3076 9824
rect 3012 9764 3016 9820
rect 3016 9764 3072 9820
rect 3072 9764 3076 9820
rect 3012 9760 3076 9764
rect 3092 9820 3156 9824
rect 3092 9764 3096 9820
rect 3096 9764 3152 9820
rect 3152 9764 3156 9820
rect 3092 9760 3156 9764
rect 3172 9820 3236 9824
rect 3172 9764 3176 9820
rect 3176 9764 3232 9820
rect 3232 9764 3236 9820
rect 3172 9760 3236 9764
rect 3252 9820 3316 9824
rect 3252 9764 3256 9820
rect 3256 9764 3312 9820
rect 3312 9764 3316 9820
rect 3252 9760 3316 9764
rect 2352 9276 2416 9280
rect 2352 9220 2356 9276
rect 2356 9220 2412 9276
rect 2412 9220 2416 9276
rect 2352 9216 2416 9220
rect 2432 9276 2496 9280
rect 2432 9220 2436 9276
rect 2436 9220 2492 9276
rect 2492 9220 2496 9276
rect 2432 9216 2496 9220
rect 2512 9276 2576 9280
rect 2512 9220 2516 9276
rect 2516 9220 2572 9276
rect 2572 9220 2576 9276
rect 2512 9216 2576 9220
rect 2592 9276 2656 9280
rect 2592 9220 2596 9276
rect 2596 9220 2652 9276
rect 2652 9220 2656 9276
rect 2592 9216 2656 9220
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 2352 8188 2416 8192
rect 2352 8132 2356 8188
rect 2356 8132 2412 8188
rect 2412 8132 2416 8188
rect 2352 8128 2416 8132
rect 2432 8188 2496 8192
rect 2432 8132 2436 8188
rect 2436 8132 2492 8188
rect 2492 8132 2496 8188
rect 2432 8128 2496 8132
rect 2512 8188 2576 8192
rect 2512 8132 2516 8188
rect 2516 8132 2572 8188
rect 2572 8132 2576 8188
rect 2512 8128 2576 8132
rect 2592 8188 2656 8192
rect 2592 8132 2596 8188
rect 2596 8132 2652 8188
rect 2652 8132 2656 8188
rect 2592 8128 2656 8132
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 2352 7100 2416 7104
rect 2352 7044 2356 7100
rect 2356 7044 2412 7100
rect 2412 7044 2416 7100
rect 2352 7040 2416 7044
rect 2432 7100 2496 7104
rect 2432 7044 2436 7100
rect 2436 7044 2492 7100
rect 2492 7044 2496 7100
rect 2432 7040 2496 7044
rect 2512 7100 2576 7104
rect 2512 7044 2516 7100
rect 2516 7044 2572 7100
rect 2572 7044 2576 7100
rect 2512 7040 2576 7044
rect 2592 7100 2656 7104
rect 2592 7044 2596 7100
rect 2596 7044 2652 7100
rect 2652 7044 2656 7100
rect 2592 7040 2656 7044
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 2352 6012 2416 6016
rect 2352 5956 2356 6012
rect 2356 5956 2412 6012
rect 2412 5956 2416 6012
rect 2352 5952 2416 5956
rect 2432 6012 2496 6016
rect 2432 5956 2436 6012
rect 2436 5956 2492 6012
rect 2492 5956 2496 6012
rect 2432 5952 2496 5956
rect 2512 6012 2576 6016
rect 2512 5956 2516 6012
rect 2516 5956 2572 6012
rect 2572 5956 2576 6012
rect 2512 5952 2576 5956
rect 2592 6012 2656 6016
rect 2592 5956 2596 6012
rect 2596 5956 2652 6012
rect 2652 5956 2656 6012
rect 2592 5952 2656 5956
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 2352 4924 2416 4928
rect 2352 4868 2356 4924
rect 2356 4868 2412 4924
rect 2412 4868 2416 4924
rect 2352 4864 2416 4868
rect 2432 4924 2496 4928
rect 2432 4868 2436 4924
rect 2436 4868 2492 4924
rect 2492 4868 2496 4924
rect 2432 4864 2496 4868
rect 2512 4924 2576 4928
rect 2512 4868 2516 4924
rect 2516 4868 2572 4924
rect 2572 4868 2576 4924
rect 2512 4864 2576 4868
rect 2592 4924 2656 4928
rect 2592 4868 2596 4924
rect 2596 4868 2652 4924
rect 2652 4868 2656 4924
rect 2592 4864 2656 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 2352 3836 2416 3840
rect 2352 3780 2356 3836
rect 2356 3780 2412 3836
rect 2412 3780 2416 3836
rect 2352 3776 2416 3780
rect 2432 3836 2496 3840
rect 2432 3780 2436 3836
rect 2436 3780 2492 3836
rect 2492 3780 2496 3836
rect 2432 3776 2496 3780
rect 2512 3836 2576 3840
rect 2512 3780 2516 3836
rect 2516 3780 2572 3836
rect 2572 3780 2576 3836
rect 2512 3776 2576 3780
rect 2592 3836 2656 3840
rect 2592 3780 2596 3836
rect 2596 3780 2652 3836
rect 2652 3780 2656 3836
rect 2592 3776 2656 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 2352 2748 2416 2752
rect 2352 2692 2356 2748
rect 2356 2692 2412 2748
rect 2412 2692 2416 2748
rect 2352 2688 2416 2692
rect 2432 2748 2496 2752
rect 2432 2692 2436 2748
rect 2436 2692 2492 2748
rect 2492 2692 2496 2748
rect 2432 2688 2496 2692
rect 2512 2748 2576 2752
rect 2512 2692 2516 2748
rect 2516 2692 2572 2748
rect 2572 2692 2576 2748
rect 2512 2688 2576 2692
rect 2592 2748 2656 2752
rect 2592 2692 2596 2748
rect 2596 2692 2652 2748
rect 2652 2692 2656 2748
rect 2592 2688 2656 2692
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
<< metal4 >>
rect 2344 20160 2664 20176
rect 2344 20096 2352 20160
rect 2416 20096 2432 20160
rect 2496 20096 2512 20160
rect 2576 20096 2592 20160
rect 2656 20096 2664 20160
rect 2344 19072 2664 20096
rect 2344 19008 2352 19072
rect 2416 19008 2432 19072
rect 2496 19008 2512 19072
rect 2576 19008 2592 19072
rect 2656 19008 2664 19072
rect 2344 17984 2664 19008
rect 2344 17920 2352 17984
rect 2416 17920 2432 17984
rect 2496 17920 2512 17984
rect 2576 17920 2592 17984
rect 2656 17920 2664 17984
rect 2344 16896 2664 17920
rect 2344 16832 2352 16896
rect 2416 16832 2432 16896
rect 2496 16832 2512 16896
rect 2576 16832 2592 16896
rect 2656 16832 2664 16896
rect 2344 15808 2664 16832
rect 2344 15744 2352 15808
rect 2416 15744 2432 15808
rect 2496 15744 2512 15808
rect 2576 15744 2592 15808
rect 2656 15744 2664 15808
rect 2344 14720 2664 15744
rect 2344 14656 2352 14720
rect 2416 14656 2432 14720
rect 2496 14656 2512 14720
rect 2576 14656 2592 14720
rect 2656 14656 2664 14720
rect 2344 13632 2664 14656
rect 2344 13568 2352 13632
rect 2416 13568 2432 13632
rect 2496 13568 2512 13632
rect 2576 13568 2592 13632
rect 2656 13568 2664 13632
rect 2344 12544 2664 13568
rect 2344 12480 2352 12544
rect 2416 12480 2432 12544
rect 2496 12480 2512 12544
rect 2576 12480 2592 12544
rect 2656 12480 2664 12544
rect 2344 11456 2664 12480
rect 2344 11392 2352 11456
rect 2416 11392 2432 11456
rect 2496 11392 2512 11456
rect 2576 11392 2592 11456
rect 2656 11392 2664 11456
rect 2344 10368 2664 11392
rect 2344 10304 2352 10368
rect 2416 10304 2432 10368
rect 2496 10304 2512 10368
rect 2576 10304 2592 10368
rect 2656 10304 2664 10368
rect 2344 9280 2664 10304
rect 2344 9216 2352 9280
rect 2416 9216 2432 9280
rect 2496 9216 2512 9280
rect 2576 9216 2592 9280
rect 2656 9216 2664 9280
rect 2344 8192 2664 9216
rect 2344 8128 2352 8192
rect 2416 8128 2432 8192
rect 2496 8128 2512 8192
rect 2576 8128 2592 8192
rect 2656 8128 2664 8192
rect 2344 7104 2664 8128
rect 2344 7040 2352 7104
rect 2416 7040 2432 7104
rect 2496 7040 2512 7104
rect 2576 7040 2592 7104
rect 2656 7040 2664 7104
rect 2344 6016 2664 7040
rect 2344 5952 2352 6016
rect 2416 5952 2432 6016
rect 2496 5952 2512 6016
rect 2576 5952 2592 6016
rect 2656 5952 2664 6016
rect 2344 4928 2664 5952
rect 2344 4864 2352 4928
rect 2416 4864 2432 4928
rect 2496 4864 2512 4928
rect 2576 4864 2592 4928
rect 2656 4864 2664 4928
rect 2344 3840 2664 4864
rect 2344 3776 2352 3840
rect 2416 3776 2432 3840
rect 2496 3776 2512 3840
rect 2576 3776 2592 3840
rect 2656 3776 2664 3840
rect 2344 3694 2664 3776
rect 2344 3458 2386 3694
rect 2622 3458 2664 3694
rect 2344 2752 2664 3458
rect 2344 2688 2352 2752
rect 2416 2688 2432 2752
rect 2496 2688 2512 2752
rect 2576 2688 2592 2752
rect 2656 2688 2664 2752
rect 2344 2128 2664 2688
rect 3004 19616 3324 20176
rect 3004 19552 3012 19616
rect 3076 19552 3092 19616
rect 3156 19552 3172 19616
rect 3236 19552 3252 19616
rect 3316 19552 3324 19616
rect 3004 18528 3324 19552
rect 3004 18464 3012 18528
rect 3076 18464 3092 18528
rect 3156 18464 3172 18528
rect 3236 18464 3252 18528
rect 3316 18464 3324 18528
rect 3004 17440 3324 18464
rect 3004 17376 3012 17440
rect 3076 17376 3092 17440
rect 3156 17376 3172 17440
rect 3236 17376 3252 17440
rect 3316 17376 3324 17440
rect 3004 16352 3324 17376
rect 3004 16288 3012 16352
rect 3076 16288 3092 16352
rect 3156 16288 3172 16352
rect 3236 16288 3252 16352
rect 3316 16288 3324 16352
rect 3004 15264 3324 16288
rect 3004 15200 3012 15264
rect 3076 15200 3092 15264
rect 3156 15200 3172 15264
rect 3236 15200 3252 15264
rect 3316 15200 3324 15264
rect 3004 14176 3324 15200
rect 3004 14112 3012 14176
rect 3076 14112 3092 14176
rect 3156 14112 3172 14176
rect 3236 14112 3252 14176
rect 3316 14112 3324 14176
rect 3004 13088 3324 14112
rect 3004 13024 3012 13088
rect 3076 13024 3092 13088
rect 3156 13024 3172 13088
rect 3236 13024 3252 13088
rect 3316 13024 3324 13088
rect 3004 12000 3324 13024
rect 3004 11936 3012 12000
rect 3076 11936 3092 12000
rect 3156 11936 3172 12000
rect 3236 11936 3252 12000
rect 3316 11936 3324 12000
rect 3004 10912 3324 11936
rect 3004 10848 3012 10912
rect 3076 10848 3092 10912
rect 3156 10848 3172 10912
rect 3236 10848 3252 10912
rect 3316 10848 3324 10912
rect 3004 9824 3324 10848
rect 3004 9760 3012 9824
rect 3076 9760 3092 9824
rect 3156 9760 3172 9824
rect 3236 9760 3252 9824
rect 3316 9760 3324 9824
rect 3004 8736 3324 9760
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4354 3092 4384
rect 3156 4354 3172 4384
rect 3236 4354 3252 4384
rect 3316 4320 3324 4384
rect 3004 4118 3046 4320
rect 3282 4118 3324 4320
rect 3004 3296 3324 4118
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 2128 3324 2144
<< via4 >>
rect 2386 3458 2622 3694
rect 3046 4320 3076 4354
rect 3076 4320 3092 4354
rect 3092 4320 3156 4354
rect 3156 4320 3172 4354
rect 3172 4320 3236 4354
rect 3236 4320 3252 4354
rect 3252 4320 3282 4354
rect 3046 4118 3282 4320
<< metal5 >>
rect 1056 4354 19184 4396
rect 1056 4118 3046 4354
rect 3282 4118 19184 4354
rect 1056 4076 19184 4118
rect 1056 3694 19184 3736
rect 1056 3458 2386 3694
rect 2622 3458 19184 3694
rect 1056 3416 19184 3458
use sky130_fd_sc_hd__inv_2  _194_
timestamp -3599
transform 1 0 4968 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _195_
timestamp -3599
transform 1 0 11684 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _196_
timestamp -3599
transform -1 0 3680 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _197_
timestamp -3599
transform -1 0 4876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _198_
timestamp -3599
transform -1 0 4692 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _199_
timestamp -3599
transform 1 0 2760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _200_
timestamp -3599
transform 1 0 3496 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _201_
timestamp -3599
transform -1 0 7452 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _202_
timestamp -3599
transform -1 0 11776 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _203_
timestamp -3599
transform 1 0 10120 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _204_
timestamp -3599
transform 1 0 10396 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _205_
timestamp -3599
transform -1 0 13064 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _206_
timestamp -3599
transform 1 0 12144 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _207_
timestamp -3599
transform -1 0 16192 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _208_
timestamp -3599
transform 1 0 15088 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _209_
timestamp -3599
transform 1 0 14996 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _210_
timestamp -3599
transform -1 0 18308 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _211_
timestamp -3599
transform 1 0 17204 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _212_
timestamp -3599
transform -1 0 14628 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _213_
timestamp -3599
transform 1 0 16008 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _214_
timestamp -3599
transform 1 0 14076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _215_
timestamp -3599
transform -1 0 18124 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _216_
timestamp -3599
transform 1 0 17020 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _217_
timestamp -3599
transform 1 0 7176 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _218_
timestamp -3599
transform 1 0 6532 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _219_
timestamp -3599
transform 1 0 7176 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _220_
timestamp -3599
transform -1 0 9384 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _221_
timestamp -3599
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _222_
timestamp -3599
transform -1 0 15456 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _223_
timestamp -3599
transform 1 0 14536 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _224_
timestamp -3599
transform 1 0 14628 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _225_
timestamp -3599
transform -1 0 16836 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _226_
timestamp -3599
transform -1 0 17020 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _227_
timestamp -3599
transform -1 0 9108 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _228_
timestamp -3599
transform -1 0 8832 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _229_
timestamp -3599
transform -1 0 14720 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _230_
timestamp -3599
transform 1 0 16652 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _231_
timestamp -3599
transform 1 0 13432 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _232_
timestamp -3599
transform -1 0 18308 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _233_
timestamp -3599
transform 1 0 17112 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _234_
timestamp -3599
transform 1 0 5704 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _235_
timestamp -3599
transform -1 0 6992 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _236_
timestamp -3599
transform 1 0 5520 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _237_
timestamp -3599
transform -1 0 8464 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _238_
timestamp -3599
transform -1 0 8004 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _239_
timestamp -3599
transform 1 0 8372 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _240_
timestamp -3599
transform -1 0 8832 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _241_
timestamp -3599
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _242_
timestamp -3599
transform -1 0 9844 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _243_
timestamp -3599
transform -1 0 9660 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _244_
timestamp -3599
transform -1 0 14352 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _245_
timestamp -3599
transform 1 0 16744 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _246_
timestamp -3599
transform 1 0 14076 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _247_
timestamp -3599
transform -1 0 18400 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _248_
timestamp -3599
transform 1 0 17204 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _249_
timestamp -3599
transform -1 0 3128 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _250_
timestamp -3599
transform -1 0 2208 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _251_
timestamp -3599
transform 1 0 2300 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _252_
timestamp -3599
transform 1 0 2024 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _253_
timestamp -3599
transform 1 0 2024 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _254_
timestamp -3599
transform 1 0 15272 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _255_
timestamp -3599
transform 1 0 16192 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _256_
timestamp -3599
transform 1 0 15180 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _257_
timestamp -3599
transform -1 0 18216 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _258_
timestamp -3599
transform 1 0 17112 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _259_
timestamp -3599
transform -1 0 11500 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _260_
timestamp -3599
transform 1 0 10488 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _261_
timestamp -3599
transform -1 0 11224 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _262_
timestamp -3599
transform -1 0 12144 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _263_
timestamp -3599
transform 1 0 12236 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _264_
timestamp -3599
transform -1 0 15456 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _265_
timestamp -3599
transform 1 0 15456 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _266_
timestamp -3599
transform 1 0 14628 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _267_
timestamp -3599
transform -1 0 18216 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _268_
timestamp -3599
transform 1 0 17020 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _269_
timestamp -3599
transform -1 0 4416 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _270_
timestamp -3599
transform 1 0 4324 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _271_
timestamp -3599
transform -1 0 3772 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _272_
timestamp -3599
transform -1 0 2392 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _273_
timestamp -3599
transform 1 0 3772 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _274_
timestamp -3599
transform -1 0 7636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _275_
timestamp -3599
transform 1 0 6440 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _276_
timestamp -3599
transform 1 0 6440 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _277_
timestamp -3599
transform 1 0 2760 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _278_
timestamp -3599
transform -1 0 4968 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _279_
timestamp -3599
transform -1 0 4416 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _280_
timestamp -3599
transform 1 0 4416 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_1  _281_
timestamp -3599
transform 1 0 4968 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _282_
timestamp -3599
transform -1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _283_
timestamp -3599
transform 1 0 1472 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _284_
timestamp -3599
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _285_
timestamp -3599
transform 1 0 3772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _286_
timestamp -3599
transform -1 0 3496 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _287_
timestamp -3599
transform 1 0 6348 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _288_
timestamp -3599
transform 1 0 2944 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _289_
timestamp -3599
transform 1 0 3772 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _290_
timestamp -3599
transform 1 0 4048 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _291_
timestamp -3599
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_1  _292_
timestamp -3599
transform -1 0 4232 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _293_
timestamp -3599
transform 1 0 6348 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _294_
timestamp -3599
transform 1 0 15916 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _295_
timestamp -3599
transform -1 0 12328 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _296_
timestamp -3599
transform 1 0 16192 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _297_
timestamp -3599
transform 1 0 14628 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _298_
timestamp -3599
transform 1 0 7268 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _299_
timestamp -3599
transform 1 0 15088 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _300_
timestamp -3599
transform 1 0 15272 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _301_
timestamp -3599
transform 1 0 6348 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _302_
timestamp -3599
transform 1 0 9016 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _303_
timestamp -3599
transform 1 0 14904 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _304_
timestamp -3599
transform -1 0 4692 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _305_
timestamp -3599
transform 1 0 15364 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _306_
timestamp -3599
transform -1 0 12512 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _307_
timestamp -3599
transform 1 0 8924 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _308_
timestamp -3599
transform 1 0 4968 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _309_
timestamp -3599
transform 1 0 4784 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _310_
timestamp -3599
transform -1 0 2116 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _311_
timestamp -3599
transform 1 0 3312 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _312_
timestamp -3599
transform 1 0 1932 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _313_
timestamp -3599
transform 1 0 3312 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _314_
timestamp -3599
transform 1 0 3772 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _315_
timestamp -3599
transform 1 0 2576 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _316_
timestamp -3599
transform 1 0 3680 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp -3599
transform -1 0 13156 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _318_
timestamp -3599
transform -1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp -3599
transform -1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp -3599
transform -1 0 6164 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp -3599
transform 1 0 2484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp -3599
transform 1 0 2300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp -3599
transform -1 0 5612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp -3599
transform 1 0 2852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp -3599
transform 1 0 2300 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp -3599
transform -1 0 7636 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp -3599
transform -1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp -3599
transform 1 0 2392 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp -3599
transform -1 0 6440 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp -3599
transform -1 0 3220 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _331_
timestamp -3599
transform -1 0 5612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp -3599
transform -1 0 2300 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp -3599
transform -1 0 5520 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp -3599
transform -1 0 7268 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp -3599
transform -1 0 11132 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp -3599
transform 1 0 8464 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp -3599
transform -1 0 5888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp -3599
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp -3599
transform 1 0 12512 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp -3599
transform -1 0 18492 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp -3599
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp -3599
transform 1 0 18400 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp -3599
transform 1 0 14996 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp -3599
transform -1 0 13524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp -3599
transform -1 0 11132 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp -3599
transform -1 0 4048 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp -3599
transform 1 0 3956 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp -3599
transform 1 0 17940 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp -3599
transform -1 0 15824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp -3599
transform 1 0 17388 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp -3599
transform 1 0 14444 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp -3599
transform 1 0 2668 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp -3599
transform -1 0 3404 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp -3599
transform -1 0 9752 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _355_
timestamp -3599
transform -1 0 9200 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp -3599
transform 1 0 18400 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp -3599
transform 1 0 13248 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp -3599
transform 1 0 7176 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp -3599
transform -1 0 6256 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp -3599
transform -1 0 11776 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _361_
timestamp -3599
transform -1 0 9660 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp -3599
transform -1 0 18400 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp -3599
transform -1 0 16192 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp -3599
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp -3599
transform -1 0 5704 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp -3599
transform 1 0 16836 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _367_
timestamp -3599
transform -1 0 14904 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp -3599
transform 1 0 17940 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp -3599
transform -1 0 14352 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _370_
timestamp -3599
transform 1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp -3599
transform 1 0 8096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp -3599
transform 1 0 6992 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _373_
timestamp -3599
transform 1 0 17572 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp -3599
transform -1 0 15456 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp -3599
transform 1 0 17204 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _376_
timestamp -3599
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _377_
timestamp -3599
transform -1 0 9936 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _378_
timestamp -3599
transform -1 0 8372 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _379_
timestamp -3599
transform 1 0 17204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _380_
timestamp -3599
transform 1 0 15364 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _381_
timestamp -3599
transform 1 0 17848 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _382_
timestamp -3599
transform -1 0 14904 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _383_
timestamp -3599
transform -1 0 11776 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _384_
timestamp -3599
transform -1 0 12788 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _385_
timestamp -3599
transform 1 0 18400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _386_
timestamp -3599
transform -1 0 16008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _387_
timestamp -3599
transform -1 0 16928 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _388_
timestamp -3599
transform -1 0 16284 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _389_
timestamp -3599
transform 1 0 12972 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _390_
timestamp -3599
transform -1 0 11224 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _391_
timestamp -3599
transform 1 0 5520 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _392_
timestamp -3599
transform -1 0 13984 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _393_
timestamp -3599
transform -1 0 3220 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _394_
timestamp -3599
transform 1 0 3680 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _395_
timestamp -3599
transform 1 0 4048 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _396_
timestamp -3599
transform 1 0 1472 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _397_
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _398_
timestamp -3599
transform 1 0 4232 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _399_
timestamp -3599
transform 1 0 1840 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _400_
timestamp -3599
transform 1 0 1380 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _401_
timestamp -3599
transform 1 0 5520 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _402_
timestamp -3599
transform 1 0 3864 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _403_
timestamp -3599
transform 1 0 1380 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _404_
timestamp -3599
transform 1 0 4324 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _405_
timestamp -3599
transform 1 0 1840 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _406_
timestamp -3599
transform 1 0 3496 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _407_
timestamp -3599
transform 1 0 1380 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _408_
timestamp -3599
transform -1 0 5888 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _409_
timestamp -3599
transform 1 0 5520 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _410_
timestamp -3599
transform 1 0 9016 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _411_
timestamp -3599
transform 1 0 7452 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _412_
timestamp -3599
transform 1 0 3772 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _413_
timestamp -3599
transform 1 0 11500 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _414_
timestamp -3599
transform 1 0 11500 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _415_
timestamp -3599
transform 1 0 16836 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _416_
timestamp -3599
transform 1 0 14076 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _417_
timestamp -3599
transform 1 0 16560 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _418_
timestamp -3599
transform 1 0 14076 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _419_
timestamp -3599
transform 1 0 12144 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _420_
timestamp -3599
transform -1 0 11408 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _421_
timestamp -3599
transform 1 0 2668 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _422_
timestamp -3599
transform 1 0 3128 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _423_
timestamp -3599
transform 1 0 16928 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _424_
timestamp -3599
transform 1 0 14260 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _425_
timestamp -3599
transform 1 0 16652 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _426_
timestamp -3599
transform -1 0 16008 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _427_
timestamp -3599
transform 1 0 1656 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _428_
timestamp -3599
transform 1 0 1748 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _429_
timestamp -3599
transform 1 0 7728 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _430_
timestamp -3599
transform 1 0 7728 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _431_
timestamp -3599
transform 1 0 17020 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _432_
timestamp -3599
transform 1 0 12328 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _433_
timestamp -3599
transform 1 0 6164 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _434_
timestamp -3599
transform 1 0 4692 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _435_
timestamp -3599
transform 1 0 9660 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _436_
timestamp -3599
transform 1 0 7544 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _437_
timestamp -3599
transform 1 0 16284 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _438_
timestamp -3599
transform 1 0 14720 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _439_
timestamp -3599
transform 1 0 7544 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _440_
timestamp -3599
transform 1 0 4324 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _441_
timestamp -3599
transform 1 0 16652 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _442_
timestamp -3599
transform -1 0 15916 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _443_
timestamp -3599
transform 1 0 17020 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _444_
timestamp -3599
transform 1 0 12880 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _445_
timestamp -3599
transform 1 0 8924 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _446_
timestamp -3599
transform 1 0 7084 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _447_
timestamp -3599
transform 1 0 5980 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _448_
timestamp -3599
transform 1 0 16652 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _449_
timestamp -3599
transform 1 0 14076 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _450_
timestamp -3599
transform 1 0 16652 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _451_
timestamp -3599
transform -1 0 15916 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _452_
timestamp -3599
transform 1 0 7728 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _453_
timestamp -3599
transform 1 0 6256 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _454_
timestamp -3599
transform 1 0 16652 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _455_
timestamp -3599
transform 1 0 14352 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _456_
timestamp -3599
transform 1 0 16836 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _457_
timestamp -3599
transform 1 0 12144 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _458_
timestamp -3599
transform 1 0 9568 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _459_
timestamp -3599
transform 1 0 10672 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _460_
timestamp -3599
transform 1 0 17020 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _461_
timestamp -3599
transform 1 0 14076 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _462_
timestamp -3599
transform 1 0 15548 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _463_
timestamp -3599
transform 1 0 14168 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _464_
timestamp -3599
transform 1 0 11960 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _465_
timestamp -3599
transform 1 0 9568 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _466_
timestamp -3599
transform -1 0 10672 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _467_
timestamp -3599
transform -1 0 13984 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _468_
timestamp -3599
transform -1 0 18400 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _469_
timestamp -3599
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _470_
timestamp -3599
transform 1 0 18492 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _471_
timestamp -3599
transform -1 0 12236 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _472_
timestamp -3599
transform -1 0 9476 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _473_
timestamp -3599
transform 1 0 18124 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _474_
timestamp -3599
transform 1 0 18124 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _475_
timestamp -3599
transform -1 0 10304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _476_
timestamp -3599
transform -1 0 18676 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _477_
timestamp -3599
transform -1 0 18400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _478_
timestamp -3599
transform -1 0 13892 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _479_
timestamp -3599
transform -1 0 18400 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _480_
timestamp -3599
transform 1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _481_
timestamp -3599
transform 1 0 1564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _482_
timestamp -3599
transform 1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _483_
timestamp -3599
transform 1 0 1748 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _484_
timestamp -3599
transform -1 0 11776 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _485_
timestamp -3599
transform -1 0 13616 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _486_
timestamp -3599
transform -1 0 18400 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _487_
timestamp -3599
transform -1 0 4968 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _488_
timestamp -3599
transform 1 0 18400 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _489_
timestamp -3599
transform -1 0 11408 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _490_
timestamp -3599
transform -1 0 8280 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _491_
timestamp -3599
transform -1 0 18676 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _492_
timestamp -3599
transform -1 0 18676 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _493_
timestamp -3599
transform -1 0 9200 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _494_
timestamp -3599
transform 1 0 18492 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _495_
timestamp -3599
transform -1 0 18768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _496_
timestamp -3599
transform -1 0 13340 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _497_
timestamp -3599
transform -1 0 18400 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _498_
timestamp -3599
transform -1 0 6072 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _499_
timestamp -3599
transform 1 0 2300 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _500_
timestamp -3599
transform 1 0 5244 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _501_
timestamp -3599
transform 1 0 5428 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _502_
timestamp -3599
transform 1 0 9292 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _503_
timestamp -3599
transform 1 0 11960 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _504_
timestamp -3599
transform 1 0 15824 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _505_
timestamp -3599
transform -1 0 4140 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _506_
timestamp -3599
transform 1 0 16008 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _507_
timestamp -3599
transform 1 0 9568 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _508_
timestamp -3599
transform 1 0 6532 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _509_
timestamp -3599
transform 1 0 15456 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _510_
timestamp -3599
transform 1 0 15548 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _511_
timestamp -3599
transform 1 0 7544 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _512_
timestamp -3599
transform 1 0 14812 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _513_
timestamp -3599
transform 1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _514_
timestamp -3599
transform 1 0 11776 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _515_
timestamp -3599
transform 1 0 15548 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp -3599
transform 1 0 9292 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp -3599
transform -1 0 8188 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp -3599
transform -1 0 8188 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp -3599
transform 1 0 12512 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp -3599
transform 1 0 13156 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp -3599
transform -1 0 6900 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp -3599
transform -1 0 8372 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp -3599
transform 1 0 14076 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp -3599
transform 1 0 14168 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__bufinv_16  clkload0
timestamp -3599
transform 1 0 5520 0 1 8704
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_4  clkload1
timestamp -3599
transform -1 0 13064 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__bufinv_16  clkload2
timestamp -3599
transform 1 0 13156 0 -1 8704
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinvlp_4  clkload3
timestamp -3599
transform 1 0 5612 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  clkload4
timestamp -3599
transform 1 0 6532 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__bufinv_16  clkload5
timestamp -3599
transform 1 0 13340 0 -1 14144
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_4  clkload6
timestamp -3599
transform -1 0 13156 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636964856
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636964856
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -3599
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636964856
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41
timestamp -3599
transform 1 0 4876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49
timestamp -3599
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp -3599
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp -3599
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62
timestamp -3599
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69
timestamp -3599
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79
timestamp -3599
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp -3599
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp -3599
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_90
timestamp -3599
transform 1 0 9384 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_98
timestamp -3599
transform 1 0 10120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104
timestamp -3599
transform 1 0 10672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp -3599
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp -3599
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121
timestamp -3599
transform 1 0 12236 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_125
timestamp -3599
transform 1 0 12604 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_133
timestamp -3599
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp -3599
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp -3599
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_146
timestamp -3599
transform 1 0 14536 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_154
timestamp -3599
transform 1 0 15272 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_160
timestamp -3599
transform 1 0 15824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_169
timestamp -3599
transform 1 0 16652 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6
timestamp 1636964856
transform 1 0 1656 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_18
timestamp -3599
transform 1 0 2760 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_26
timestamp -3599
transform 1 0 3496 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp -3599
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_57
timestamp -3599
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_88
timestamp -3599
transform 1 0 9200 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_92
timestamp -3599
transform 1 0 9568 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_96
timestamp -3599
transform 1 0 9936 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_100
timestamp -3599
transform 1 0 10304 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_136
timestamp -3599
transform 1 0 13616 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_140
timestamp 1636964856
transform 1 0 13984 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_162
timestamp -3599
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_192
timestamp -3599
transform 1 0 18768 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_23
timestamp -3599
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -3599
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_32
timestamp 1636964856
transform 1 0 4048 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_44
timestamp -3599
transform 1 0 5152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_71
timestamp -3599
transform 1 0 7636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_75
timestamp -3599
transform 1 0 8004 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_105
timestamp -3599
transform 1 0 10764 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_113
timestamp -3599
transform 1 0 11500 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_164
timestamp -3599
transform 1 0 16192 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_172
timestamp -3599
transform 1 0 16928 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_183
timestamp -3599
transform 1 0 17940 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_191
timestamp -3599
transform 1 0 18676 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp -3599
transform 1 0 1380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_13
timestamp -3599
transform 1 0 2300 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_21
timestamp -3599
transform 1 0 3036 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_49
timestamp -3599
transform 1 0 5612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp -3599
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp -3599
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_67
timestamp -3599
transform 1 0 7268 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_78
timestamp -3599
transform 1 0 8280 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_87
timestamp 1636964856
transform 1 0 9108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_99
timestamp 1636964856
transform 1 0 10212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp -3599
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_113
timestamp -3599
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_129
timestamp -3599
transform 1 0 12972 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_135
timestamp 1636964856
transform 1 0 13524 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_147
timestamp -3599
transform 1 0 14628 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_157
timestamp -3599
transform 1 0 15548 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_169
timestamp -3599
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_21
timestamp -3599
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -3599
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_35
timestamp 1636964856
transform 1 0 4324 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_47
timestamp -3599
transform 1 0 5428 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_73
timestamp -3599
transform 1 0 7820 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp -3599
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_85
timestamp -3599
transform 1 0 8924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_94
timestamp -3599
transform 1 0 9752 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_102
timestamp -3599
transform 1 0 10488 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_113
timestamp -3599
transform 1 0 11500 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_117
timestamp -3599
transform 1 0 11868 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_126
timestamp 1636964856
transform 1 0 12696 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp -3599
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_141
timestamp -3599
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_169
timestamp 1636964856
transform 1 0 16652 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_181
timestamp -3599
transform 1 0 17756 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_187
timestamp -3599
transform 1 0 18308 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp -3599
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_30
timestamp -3599
transform 1 0 3864 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_38
timestamp -3599
transform 1 0 4600 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp -3599
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_57
timestamp -3599
transform 1 0 6348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_63
timestamp -3599
transform 1 0 6900 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_133
timestamp 1636964856
transform 1 0 13340 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_145
timestamp -3599
transform 1 0 14444 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_152
timestamp -3599
transform 1 0 15088 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_158
timestamp -3599
transform 1 0 15640 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp -3599
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp -3599
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_181
timestamp -3599
transform 1 0 17756 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_185
timestamp -3599
transform 1 0 18124 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_189
timestamp -3599
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_17
timestamp -3599
transform 1 0 2668 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp -3599
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_55
timestamp -3599
transform 1 0 6164 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_91
timestamp 1636964856
transform 1 0 9476 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_103
timestamp -3599
transform 1 0 10580 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_109
timestamp -3599
transform 1 0 11132 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_117
timestamp -3599
transform 1 0 11868 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_127
timestamp -3599
transform 1 0 12788 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_135
timestamp -3599
transform 1 0 13524 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_161
timestamp -3599
transform 1 0 15916 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_169
timestamp -3599
transform 1 0 16652 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_191
timestamp -3599
transform 1 0 18676 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_10
timestamp -3599
transform 1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_16
timestamp -3599
transform 1 0 2576 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_26
timestamp 1636964856
transform 1 0 3496 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_38
timestamp 1636964856
transform 1 0 4600 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp -3599
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636964856
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_69
timestamp -3599
transform 1 0 7452 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1636964856
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp -3599
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp -3599
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_113
timestamp -3599
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_121
timestamp -3599
transform 1 0 12236 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_147
timestamp -3599
transform 1 0 14628 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_157
timestamp -3599
transform 1 0 15548 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp -3599
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_172
timestamp -3599
transform 1 0 16928 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_185
timestamp -3599
transform 1 0 18124 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_189
timestamp -3599
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp -3599
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp -3599
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_35
timestamp 1636964856
transform 1 0 4324 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_47
timestamp -3599
transform 1 0 5428 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_68
timestamp -3599
transform 1 0 7360 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_76
timestamp -3599
transform 1 0 8096 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp -3599
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_85
timestamp -3599
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_91
timestamp 1636964856
transform 1 0 9476 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_103
timestamp 1636964856
transform 1 0 10580 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_115
timestamp -3599
transform 1 0 11684 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_119
timestamp -3599
transform 1 0 12052 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_150
timestamp -3599
transform 1 0 14904 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_156
timestamp -3599
transform 1 0 15456 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_177
timestamp -3599
transform 1 0 17388 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_191
timestamp -3599
transform 1 0 18676 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6
timestamp 1636964856
transform 1 0 1656 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_18
timestamp -3599
transform 1 0 2760 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_41
timestamp -3599
transform 1 0 4876 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_45
timestamp -3599
transform 1 0 5244 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp -3599
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp -3599
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_69
timestamp -3599
transform 1 0 7452 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_100
timestamp 1636964856
transform 1 0 10304 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_113
timestamp -3599
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_121
timestamp -3599
transform 1 0 12236 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_130
timestamp 1636964856
transform 1 0 13064 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_142
timestamp -3599
transform 1 0 14168 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_146
timestamp -3599
transform 1 0 14536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp -3599
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp -3599
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1636964856
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_181
timestamp -3599
transform 1 0 17756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp -3599
transform 1 0 18400 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_11
timestamp -3599
transform 1 0 2116 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_18
timestamp -3599
transform 1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp -3599
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_54
timestamp 1636964856
transform 1 0 6072 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_66
timestamp 1636964856
transform 1 0 7176 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_78
timestamp -3599
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_88
timestamp 1636964856
transform 1 0 9200 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_100
timestamp 1636964856
transform 1 0 10304 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_112
timestamp 1636964856
transform 1 0 11408 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_124
timestamp 1636964856
transform 1 0 12512 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_136
timestamp -3599
transform 1 0 13616 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_166
timestamp -3599
transform 1 0 16376 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_172
timestamp -3599
transform 1 0 16928 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_189
timestamp -3599
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_23
timestamp -3599
transform 1 0 3220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_35
timestamp -3599
transform 1 0 4324 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1636964856
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp -3599
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp -3599
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_77
timestamp 1636964856
transform 1 0 8188 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_89
timestamp -3599
transform 1 0 9292 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_95
timestamp 1636964856
transform 1 0 9844 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp -3599
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp -3599
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1636964856
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_125
timestamp -3599
transform 1 0 12604 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_155
timestamp -3599
transform 1 0 15364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_165
timestamp -3599
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp -3599
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_191
timestamp -3599
transform 1 0 18676 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_6
timestamp -3599
transform 1 0 1656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_10
timestamp -3599
transform 1 0 2024 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_18
timestamp -3599
transform 1 0 2760 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_22
timestamp -3599
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636964856
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_41
timestamp -3599
transform 1 0 4876 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_47
timestamp -3599
transform 1 0 5428 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_72
timestamp 1636964856
transform 1 0 7728 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_116
timestamp 1636964856
transform 1 0 11776 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_128
timestamp 1636964856
transform 1 0 12880 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp -3599
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_165
timestamp -3599
transform 1 0 16284 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_173
timestamp -3599
transform 1 0 17020 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_178
timestamp -3599
transform 1 0 17480 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_186
timestamp -3599
transform 1 0 18216 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_6
timestamp -3599
transform 1 0 1656 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_28
timestamp -3599
transform 1 0 3680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp -3599
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1636964856
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1636964856
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1636964856
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1636964856
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp -3599
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp -3599
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp -3599
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_117
timestamp -3599
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_121
timestamp -3599
transform 1 0 12236 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_129
timestamp -3599
transform 1 0 12972 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_151
timestamp 1636964856
transform 1 0 14996 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_163
timestamp -3599
transform 1 0 16100 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp -3599
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_192
timestamp -3599
transform 1 0 18768 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_16
timestamp 1636964856
transform 1 0 2576 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636964856
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1636964856
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1636964856
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1636964856
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp -3599
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp -3599
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1636964856
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1636964856
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1636964856
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1636964856
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp -3599
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp -3599
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1636964856
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_159
timestamp -3599
transform 1 0 15732 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_167
timestamp -3599
transform 1 0 16468 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_191
timestamp -3599
transform 1 0 18676 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_23
timestamp -3599
transform 1 0 3220 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_31
timestamp -3599
transform 1 0 3956 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp -3599
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_66
timestamp 1636964856
transform 1 0 7176 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_78
timestamp 1636964856
transform 1 0 8280 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_90
timestamp 1636964856
transform 1 0 9384 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_102
timestamp -3599
transform 1 0 10488 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp -3599
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1636964856
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1636964856
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_137
timestamp -3599
transform 1 0 13708 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_163
timestamp -3599
transform 1 0 16100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp -3599
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1636964856
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_181
timestamp -3599
transform 1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_188
timestamp -3599
transform 1 0 18400 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_6
timestamp -3599
transform 1 0 1656 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_13
timestamp -3599
transform 1 0 2300 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_17
timestamp -3599
transform 1 0 2668 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_24
timestamp -3599
transform 1 0 3312 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_29
timestamp -3599
transform 1 0 3772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_47
timestamp -3599
transform 1 0 5428 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_71
timestamp 1636964856
transform 1 0 7636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp -3599
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1636964856
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1636964856
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1636964856
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1636964856
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp -3599
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp -3599
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1636964856
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_153
timestamp -3599
transform 1 0 15180 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_160
timestamp -3599
transform 1 0 15824 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_171
timestamp -3599
transform 1 0 16836 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_182
timestamp -3599
transform 1 0 17848 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_186
timestamp -3599
transform 1 0 18216 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_23
timestamp -3599
transform 1 0 3220 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_27
timestamp -3599
transform 1 0 3588 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_48
timestamp -3599
transform 1 0 5520 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1636964856
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1636964856
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_81
timestamp -3599
transform 1 0 8556 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp -3599
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1636964856
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_125
timestamp -3599
transform 1 0 12604 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_131
timestamp 1636964856
transform 1 0 13156 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_143
timestamp -3599
transform 1 0 14260 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_154
timestamp -3599
transform 1 0 15272 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp -3599
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_192
timestamp -3599
transform 1 0 18768 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636964856
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636964856
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp -3599
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1636964856
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1636964856
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1636964856
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1636964856
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp -3599
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp -3599
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1636964856
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1636964856
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_109
timestamp -3599
transform 1 0 11132 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_161
timestamp 1636964856
transform 1 0 15916 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_173
timestamp -3599
transform 1 0 17020 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_186
timestamp -3599
transform 1 0 18216 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_9
timestamp -3599
transform 1 0 1932 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_15
timestamp -3599
transform 1 0 2484 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_24
timestamp 1636964856
transform 1 0 3312 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_36
timestamp 1636964856
transform 1 0 4416 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_48
timestamp -3599
transform 1 0 5520 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1636964856
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1636964856
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1636964856
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1636964856
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp -3599
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp -3599
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1636964856
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_125
timestamp -3599
transform 1 0 12604 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_148
timestamp -3599
transform 1 0 14720 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_159
timestamp -3599
transform 1 0 15732 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp -3599
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1636964856
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_181
timestamp -3599
transform 1 0 17756 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_188
timestamp -3599
transform 1 0 18400 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp -3599
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_58
timestamp 1636964856
transform 1 0 6440 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_70
timestamp 1636964856
transform 1 0 7544 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp -3599
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1636964856
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1636964856
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1636964856
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1636964856
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_133
timestamp -3599
transform 1 0 13340 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_164
timestamp -3599
transform 1 0 16192 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_191
timestamp -3599
transform 1 0 18676 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_10
timestamp -3599
transform 1 0 2024 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_18
timestamp -3599
transform 1 0 2760 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_23
timestamp -3599
transform 1 0 3220 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_29
timestamp -3599
transform 1 0 3772 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_36
timestamp -3599
transform 1 0 4416 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1636964856
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1636964856
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1636964856
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1636964856
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp -3599
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp -3599
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1636964856
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_125
timestamp -3599
transform 1 0 12604 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_157
timestamp -3599
transform 1 0 15548 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp -3599
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_176
timestamp -3599
transform 1 0 17296 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp -3599
transform 1 0 17848 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_186
timestamp -3599
transform 1 0 18216 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp -3599
transform 1 0 1380 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_17
timestamp -3599
transform 1 0 2668 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_25
timestamp -3599
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_38
timestamp -3599
transform 1 0 4600 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_42
timestamp -3599
transform 1 0 4968 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_63
timestamp 1636964856
transform 1 0 6900 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_75
timestamp -3599
transform 1 0 8004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp -3599
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1636964856
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1636964856
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1636964856
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1636964856
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp -3599
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp -3599
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_144
timestamp -3599
transform 1 0 14352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_168
timestamp -3599
transform 1 0 16560 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_172
timestamp -3599
transform 1 0 16928 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_23
timestamp -3599
transform 1 0 3220 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp -3599
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp -3599
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_72
timestamp 1636964856
transform 1 0 7728 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_84
timestamp 1636964856
transform 1 0 8832 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_96
timestamp 1636964856
transform 1 0 9936 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp -3599
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp -3599
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_124
timestamp 1636964856
transform 1 0 12512 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_136
timestamp -3599
transform 1 0 13616 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_140
timestamp -3599
transform 1 0 13984 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_147
timestamp -3599
transform 1 0 14628 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_155
timestamp -3599
transform 1 0 15364 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp -3599
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp -3599
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_173
timestamp -3599
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_187
timestamp -3599
transform 1 0 18308 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_6
timestamp -3599
transform 1 0 1656 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_12
timestamp -3599
transform 1 0 2208 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_16
timestamp 1636964856
transform 1 0 2576 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1636964856
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_41
timestamp -3599
transform 1 0 4876 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_52
timestamp -3599
transform 1 0 5888 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_79
timestamp -3599
transform 1 0 8372 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp -3599
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp -3599
transform 1 0 8924 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1636964856
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_121
timestamp -3599
transform 1 0 12236 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_131
timestamp -3599
transform 1 0 13156 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp -3599
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp -3599
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_141
timestamp -3599
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_180
timestamp -3599
transform 1 0 17664 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_188
timestamp -3599
transform 1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_6
timestamp -3599
transform 1 0 1656 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_15
timestamp -3599
transform 1 0 2484 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_20
timestamp -3599
transform 1 0 2944 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_42
timestamp 1636964856
transform 1 0 4968 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp -3599
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_57
timestamp -3599
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_65
timestamp -3599
transform 1 0 7084 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_97
timestamp 1636964856
transform 1 0 10028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_109
timestamp -3599
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_113
timestamp -3599
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp -3599
transform 1 0 12236 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_162
timestamp -3599
transform 1 0 16008 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_189
timestamp -3599
transform 1 0 18492 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp -3599
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp -3599
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_79
timestamp -3599
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp -3599
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_90
timestamp 1636964856
transform 1 0 9384 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_102
timestamp -3599
transform 1 0 10488 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_127
timestamp 1636964856
transform 1 0 12788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp -3599
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_144
timestamp -3599
transform 1 0 14352 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_148
timestamp -3599
transform 1 0 14720 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_155
timestamp 1636964856
transform 1 0 15364 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_167
timestamp -3599
transform 1 0 16468 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_6
timestamp -3599
transform 1 0 1656 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_18
timestamp -3599
transform 1 0 2760 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_24
timestamp -3599
transform 1 0 3312 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_33
timestamp 1636964856
transform 1 0 4140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_45
timestamp -3599
transform 1 0 5244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp -3599
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_90
timestamp -3599
transform 1 0 9384 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_116
timestamp -3599
transform 1 0 11776 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_122
timestamp 1636964856
transform 1 0 12328 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_134
timestamp 1636964856
transform 1 0 13432 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_146
timestamp -3599
transform 1 0 14536 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_150
timestamp -3599
transform 1 0 14904 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_157
timestamp -3599
transform 1 0 15548 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp -3599
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_169
timestamp -3599
transform 1 0 16652 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_191
timestamp -3599
transform 1 0 18676 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_6
timestamp 1636964856
transform 1 0 1656 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_18
timestamp -3599
transform 1 0 2760 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp -3599
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1636964856
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1636964856
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_53
timestamp -3599
transform 1 0 5980 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_62
timestamp 1636964856
transform 1 0 6808 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_74
timestamp -3599
transform 1 0 7912 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_80
timestamp -3599
transform 1 0 8464 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1636964856
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_97
timestamp -3599
transform 1 0 10028 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_110
timestamp -3599
transform 1 0 11224 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_124
timestamp 1636964856
transform 1 0 12512 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp -3599
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_161
timestamp -3599
transform 1 0 15916 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_173
timestamp -3599
transform 1 0 17020 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_182
timestamp -3599
transform 1 0 17848 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp -3599
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_12
timestamp -3599
transform 1 0 2208 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_25
timestamp 1636964856
transform 1 0 3404 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_37
timestamp -3599
transform 1 0 4508 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_45
timestamp -3599
transform 1 0 5244 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp -3599
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp -3599
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_80
timestamp -3599
transform 1 0 8464 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_91
timestamp 1636964856
transform 1 0 9476 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_103
timestamp -3599
transform 1 0 10580 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp -3599
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_113
timestamp -3599
transform 1 0 11500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_119
timestamp -3599
transform 1 0 12052 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_128
timestamp -3599
transform 1 0 12880 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_132
timestamp 1636964856
transform 1 0 13248 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_144
timestamp -3599
transform 1 0 14352 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_156
timestamp -3599
transform 1 0 15456 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_165
timestamp -3599
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_189
timestamp -3599
transform 1 0 18492 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_6
timestamp -3599
transform 1 0 1656 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp -3599
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_32
timestamp -3599
transform 1 0 4048 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_78
timestamp -3599
transform 1 0 8280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_96
timestamp -3599
transform 1 0 9936 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_105
timestamp -3599
transform 1 0 10764 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_116
timestamp -3599
transform 1 0 11776 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp -3599
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_161
timestamp -3599
transform 1 0 15916 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_165
timestamp -3599
transform 1 0 16284 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_174
timestamp -3599
transform 1 0 17112 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_191
timestamp -3599
transform 1 0 18676 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1636964856
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_15
timestamp -3599
transform 1 0 2484 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_37
timestamp -3599
transform 1 0 4508 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_42
timestamp -3599
transform 1 0 4968 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_46
timestamp -3599
transform 1 0 5336 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp -3599
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_64
timestamp -3599
transform 1 0 6992 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_69
timestamp -3599
transform 1 0 7452 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_116
timestamp -3599
transform 1 0 11776 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_124
timestamp -3599
transform 1 0 12512 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_133
timestamp -3599
transform 1 0 13340 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_139
timestamp -3599
transform 1 0 13892 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_145
timestamp -3599
transform 1 0 14444 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_156
timestamp 1636964856
transform 1 0 15456 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_192
timestamp -3599
transform 1 0 18768 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1636964856
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1636964856
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp -3599
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1636964856
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_41
timestamp -3599
transform 1 0 4876 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_48
timestamp -3599
transform 1 0 5520 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_55
timestamp -3599
transform 1 0 6164 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_57
timestamp -3599
transform 1 0 6348 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_62
timestamp -3599
transform 1 0 6808 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_69
timestamp -3599
transform 1 0 7452 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_77
timestamp -3599
transform 1 0 8188 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp -3599
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_90
timestamp -3599
transform 1 0 9384 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_97
timestamp -3599
transform 1 0 10028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_107
timestamp -3599
transform 1 0 10948 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_111
timestamp -3599
transform 1 0 11316 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_113
timestamp -3599
transform 1 0 11500 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_118
timestamp -3599
transform 1 0 11960 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_126
timestamp -3599
transform 1 0 12696 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_132
timestamp -3599
transform 1 0 13248 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp -3599
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp -3599
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_146
timestamp -3599
transform 1 0 14536 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_153
timestamp -3599
transform 1 0 15180 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_161
timestamp -3599
transform 1 0 15916 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_167
timestamp -3599
transform 1 0 16468 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_169
timestamp -3599
transform 1 0 16652 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_175
timestamp -3599
transform 1 0 17204 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_191
timestamp -3599
transform 1 0 18676 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp -3599
transform -1 0 1932 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp -3599
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp -3599
transform 1 0 15548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp -3599
transform 1 0 10672 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp -3599
transform 1 0 17480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp -3599
transform -1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp -3599
transform 1 0 1748 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp -3599
transform 1 0 11040 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp -3599
transform 1 0 18584 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp -3599
transform -1 0 1656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp -3599
transform 1 0 18584 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp -3599
transform -1 0 8096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp -3599
transform 1 0 6532 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp -3599
transform 1 0 18584 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp -3599
transform -1 0 15180 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp -3599
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  input17
timestamp -3599
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input18
timestamp -3599
transform 1 0 7176 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp -3599
transform -1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp -3599
transform -1 0 18032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp -3599
transform -1 0 13892 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp -3599
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp -3599
transform 1 0 1748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp -3599
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp -3599
transform 1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp -3599
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp -3599
transform 1 0 1380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp -3599
transform -1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp -3599
transform 1 0 1380 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input30
timestamp -3599
transform 1 0 5888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp -3599
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp -3599
transform 1 0 16192 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp -3599
transform 1 0 5888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp -3599
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp -3599
transform -1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp -3599
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp -3599
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  input38
timestamp -3599
transform 1 0 1380 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_1  output39
timestamp -3599
transform -1 0 11316 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output40
timestamp -3599
transform 1 0 18584 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output41
timestamp -3599
transform 1 0 18584 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output42
timestamp -3599
transform -1 0 14536 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output43
timestamp -3599
transform 1 0 18584 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output44
timestamp -3599
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output45
timestamp -3599
transform -1 0 1656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output46
timestamp -3599
transform -1 0 14536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output47
timestamp -3599
transform 1 0 18584 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output48
timestamp -3599
transform -1 0 1656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output49
timestamp -3599
transform 1 0 17848 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output50
timestamp -3599
transform 1 0 18584 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output51
timestamp -3599
transform -1 0 10028 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output52
timestamp -3599
transform 1 0 17572 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output53
timestamp -3599
transform 1 0 17848 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output54
timestamp -3599
transform -1 0 10672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output55
timestamp -3599
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output56
timestamp -3599
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output57
timestamp -3599
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output58
timestamp -3599
transform -1 0 11960 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output59
timestamp -3599
transform 1 0 18308 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output60
timestamp -3599
transform 1 0 18584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output61
timestamp -3599
transform -1 0 13248 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output62
timestamp -3599
transform 1 0 18584 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output63
timestamp -3599
transform -1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output64
timestamp -3599
transform -1 0 1656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output65
timestamp -3599
transform -1 0 13892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output66
timestamp -3599
transform 1 0 18584 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output67
timestamp -3599
transform -1 0 5520 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output68
timestamp -3599
transform 1 0 17296 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output69
timestamp -3599
transform -1 0 12236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output70
timestamp -3599
transform -1 0 8740 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output71
timestamp -3599
transform 1 0 18584 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output72
timestamp -3599
transform 1 0 18584 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output73
timestamp -3599
transform -1 0 9384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_33
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 19136 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_34
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 19136 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_35
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 19136 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_36
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 19136 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_37
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 19136 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_38
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 19136 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_39
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 19136 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_40
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 19136 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_41
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 19136 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_42
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 19136 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_43
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 19136 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_44
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 19136 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_45
timestamp -3599
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -3599
transform -1 0 19136 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_46
timestamp -3599
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -3599
transform -1 0 19136 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_47
timestamp -3599
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp -3599
transform -1 0 19136 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_48
timestamp -3599
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp -3599
transform -1 0 19136 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_49
timestamp -3599
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp -3599
transform -1 0 19136 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_50
timestamp -3599
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp -3599
transform -1 0 19136 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_51
timestamp -3599
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp -3599
transform -1 0 19136 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_52
timestamp -3599
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp -3599
transform -1 0 19136 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_53
timestamp -3599
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp -3599
transform -1 0 19136 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_54
timestamp -3599
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp -3599
transform -1 0 19136 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_55
timestamp -3599
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp -3599
transform -1 0 19136 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_56
timestamp -3599
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp -3599
transform -1 0 19136 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_57
timestamp -3599
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp -3599
transform -1 0 19136 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_58
timestamp -3599
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp -3599
transform -1 0 19136 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_59
timestamp -3599
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp -3599
transform -1 0 19136 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_60
timestamp -3599
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp -3599
transform -1 0 19136 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_61
timestamp -3599
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp -3599
transform -1 0 19136 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_62
timestamp -3599
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp -3599
transform -1 0 19136 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_63
timestamp -3599
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp -3599
transform -1 0 19136 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_64
timestamp -3599
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp -3599
transform -1 0 19136 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_65
timestamp -3599
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp -3599
transform -1 0 19136 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_66
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_67
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_72
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_73
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_74
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_75
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_76
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_77
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_78
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_79
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_80
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_81
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_82
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_83
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_84
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_85
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_86
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_87
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_88
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_89
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_90
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_91
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_92
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_93
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_94
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_95
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_96
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_97
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_98
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_99
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_100
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_101
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_102
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_103
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_104
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_105
timestamp -3599
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_106
timestamp -3599
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_107
timestamp -3599
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_108
timestamp -3599
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_109
timestamp -3599
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_110
timestamp -3599
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_111
timestamp -3599
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_112
timestamp -3599
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_113
timestamp -3599
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_114
timestamp -3599
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_115
timestamp -3599
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_116
timestamp -3599
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_117
timestamp -3599
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_118
timestamp -3599
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_119
timestamp -3599
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_120
timestamp -3599
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_121
timestamp -3599
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_122
timestamp -3599
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_123
timestamp -3599
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_124
timestamp -3599
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_125
timestamp -3599
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_126
timestamp -3599
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_127
timestamp -3599
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_128
timestamp -3599
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_129
timestamp -3599
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_130
timestamp -3599
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_131
timestamp -3599
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_132
timestamp -3599
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_133
timestamp -3599
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_134
timestamp -3599
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_135
timestamp -3599
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_136
timestamp -3599
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_137
timestamp -3599
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_138
timestamp -3599
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_139
timestamp -3599
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_140
timestamp -3599
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_141
timestamp -3599
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_142
timestamp -3599
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_143
timestamp -3599
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_144
timestamp -3599
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_145
timestamp -3599
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_146
timestamp -3599
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_147
timestamp -3599
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_148
timestamp -3599
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_149
timestamp -3599
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_150
timestamp -3599
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_151
timestamp -3599
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_152
timestamp -3599
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_153
timestamp -3599
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_154
timestamp -3599
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_155
timestamp -3599
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_156
timestamp -3599
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_157
timestamp -3599
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_158
timestamp -3599
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_159
timestamp -3599
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_160
timestamp -3599
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_161
timestamp -3599
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_162
timestamp -3599
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_163
timestamp -3599
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_164
timestamp -3599
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_165
timestamp -3599
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_166
timestamp -3599
transform 1 0 6256 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_167
timestamp -3599
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_168
timestamp -3599
transform 1 0 11408 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_169
timestamp -3599
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_170
timestamp -3599
transform 1 0 16560 0 1 19584
box -38 -48 130 592
<< labels >>
flabel metal2 s 10966 21601 11022 22401 0 FreeSans 224 90 0 0 Data_in[0]
port 0 nsew signal output
flabel metal3 s 19457 7488 20257 7608 0 FreeSans 480 0 0 0 Data_in[10]
port 1 nsew signal output
flabel metal3 s 19457 4088 20257 4208 0 FreeSans 480 0 0 0 Data_in[11]
port 2 nsew signal output
flabel metal2 s 14186 21601 14242 22401 0 FreeSans 224 90 0 0 Data_in[12]
port 3 nsew signal output
flabel metal3 s 19457 5448 20257 5568 0 FreeSans 480 0 0 0 Data_in[13]
port 4 nsew signal output
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 Data_in[14]
port 5 nsew signal output
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 Data_in[15]
port 6 nsew signal output
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 Data_in[1]
port 7 nsew signal output
flabel metal3 s 19457 14968 20257 15088 0 FreeSans 480 0 0 0 Data_in[2]
port 8 nsew signal output
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 Data_in[3]
port 9 nsew signal output
flabel metal3 s 19457 19728 20257 19848 0 FreeSans 480 0 0 0 Data_in[4]
port 10 nsew signal output
flabel metal3 s 19457 10208 20257 10328 0 FreeSans 480 0 0 0 Data_in[5]
port 11 nsew signal output
flabel metal2 s 9678 21601 9734 22401 0 FreeSans 224 90 0 0 Data_in[6]
port 12 nsew signal output
flabel metal3 s 19457 21088 20257 21208 0 FreeSans 480 0 0 0 Data_in[7]
port 13 nsew signal output
flabel metal3 s 19457 19048 20257 19168 0 FreeSans 480 0 0 0 Data_in[8]
port 14 nsew signal output
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 Data_in[9]
port 15 nsew signal output
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 Data_out[0]
port 16 nsew signal input
flabel metal3 s 19457 2728 20257 2848 0 FreeSans 480 0 0 0 Data_out[10]
port 17 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 Data_out[11]
port 18 nsew signal input
flabel metal2 s 10322 21601 10378 22401 0 FreeSans 224 90 0 0 Data_out[12]
port 19 nsew signal input
flabel metal3 s 19457 1368 20257 1488 0 FreeSans 480 0 0 0 Data_out[13]
port 20 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 Data_out[14]
port 21 nsew signal input
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 Data_out[15]
port 22 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 Data_out[1]
port 23 nsew signal input
flabel metal3 s 19457 10888 20257 11008 0 FreeSans 480 0 0 0 Data_out[2]
port 24 nsew signal input
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 Data_out[3]
port 25 nsew signal input
flabel metal3 s 19457 12928 20257 13048 0 FreeSans 480 0 0 0 Data_out[4]
port 26 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 Data_out[5]
port 27 nsew signal input
flabel metal2 s 6458 21601 6514 22401 0 FreeSans 224 90 0 0 Data_out[6]
port 28 nsew signal input
flabel metal3 s 19457 14288 20257 14408 0 FreeSans 480 0 0 0 Data_out[7]
port 29 nsew signal input
flabel metal2 s 14830 21601 14886 22401 0 FreeSans 224 90 0 0 Data_out[8]
port 30 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 Data_out[9]
port 31 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 Enable
port 32 nsew signal input
flabel metal2 s 7102 21601 7158 22401 0 FreeSans 224 90 0 0 Function[0]
port 33 nsew signal input
flabel metal3 s 19457 8 20257 128 0 FreeSans 480 0 0 0 Function[10]
port 34 nsew signal input
flabel metal3 s 19457 688 20257 808 0 FreeSans 480 0 0 0 Function[11]
port 35 nsew signal input
flabel metal2 s 13542 21601 13598 22401 0 FreeSans 224 90 0 0 Function[12]
port 36 nsew signal input
flabel metal3 s 19457 6128 20257 6248 0 FreeSans 480 0 0 0 Function[13]
port 37 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 Function[14]
port 38 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 Function[15]
port 39 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 Function[1]
port 40 nsew signal input
flabel metal3 s 19457 12248 20257 12368 0 FreeSans 480 0 0 0 Function[2]
port 41 nsew signal input
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 Function[3]
port 42 nsew signal input
flabel metal3 s 19457 16328 20257 16448 0 FreeSans 480 0 0 0 Function[4]
port 43 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 Function[5]
port 44 nsew signal input
flabel metal2 s 5814 21601 5870 22401 0 FreeSans 224 90 0 0 Function[6]
port 45 nsew signal input
flabel metal3 s 19457 15648 20257 15768 0 FreeSans 480 0 0 0 Function[7]
port 46 nsew signal input
flabel metal2 s 16118 21601 16174 22401 0 FreeSans 224 90 0 0 Function[8]
port 47 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 Function[9]
port 48 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 IRQ_INT[0]
port 49 nsew signal output
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 IRQ_INT[1]
port 50 nsew signal output
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 IRQ_PIN_CHANGE
port 51 nsew signal output
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 Int_Mask[0]
port 52 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 Int_Mask[1]
port 53 nsew signal input
flabel metal2 s 9034 21601 9090 22401 0 FreeSans 224 90 0 0 PIN_DATA[0]
port 54 nsew signal bidirectional
flabel metal3 s 19457 2048 20257 2168 0 FreeSans 480 0 0 0 PIN_DATA[10]
port 55 nsew signal bidirectional
flabel metal3 s 19457 4768 20257 4888 0 FreeSans 480 0 0 0 PIN_DATA[11]
port 56 nsew signal bidirectional
flabel metal2 s 12254 21601 12310 22401 0 FreeSans 224 90 0 0 PIN_DATA[12]
port 57 nsew signal bidirectional
flabel metal3 s 19457 8168 20257 8288 0 FreeSans 480 0 0 0 PIN_DATA[13]
port 58 nsew signal bidirectional
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 PIN_DATA[14]
port 59 nsew signal bidirectional
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 PIN_DATA[15]
port 60 nsew signal bidirectional
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 PIN_DATA[1]
port 61 nsew signal bidirectional
flabel metal3 s 19457 11568 20257 11688 0 FreeSans 480 0 0 0 PIN_DATA[2]
port 62 nsew signal bidirectional
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 PIN_DATA[3]
port 63 nsew signal bidirectional
flabel metal3 s 19457 17008 20257 17128 0 FreeSans 480 0 0 0 PIN_DATA[4]
port 64 nsew signal bidirectional
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 PIN_DATA[5]
port 65 nsew signal bidirectional
flabel metal2 s 7746 21601 7802 22401 0 FreeSans 224 90 0 0 PIN_DATA[6]
port 66 nsew signal bidirectional
flabel metal3 s 19457 20408 20257 20528 0 FreeSans 480 0 0 0 PIN_DATA[7]
port 67 nsew signal bidirectional
flabel metal3 s 19457 17688 20257 17808 0 FreeSans 480 0 0 0 PIN_DATA[8]
port 68 nsew signal bidirectional
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 PIN_DATA[9]
port 69 nsew signal bidirectional
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 Pin_Change_Mask[0]
port 70 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 Pin_Change_Mask[10]
port 71 nsew signal input
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 Pin_Change_Mask[11]
port 72 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 Pin_Change_Mask[12]
port 73 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 Pin_Change_Mask[13]
port 74 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 Pin_Change_Mask[14]
port 75 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 Pin_Change_Mask[15]
port 76 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 Pin_Change_Mask[1]
port 77 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 Pin_Change_Mask[2]
port 78 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 Pin_Change_Mask[3]
port 79 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 Pin_Change_Mask[4]
port 80 nsew signal input
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 Pin_Change_Mask[5]
port 81 nsew signal input
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 Pin_Change_Mask[6]
port 82 nsew signal input
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 Pin_Change_Mask[7]
port 83 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 Pin_Change_Mask[8]
port 84 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 Pin_Change_Mask[9]
port 85 nsew signal input
flabel metal2 s 11610 21601 11666 22401 0 FreeSans 224 90 0 0 Pin_out[0]
port 86 nsew signal output
flabel metal3 s 19457 8848 20257 8968 0 FreeSans 480 0 0 0 Pin_out[10]
port 87 nsew signal output
flabel metal3 s 19457 3408 20257 3528 0 FreeSans 480 0 0 0 Pin_out[11]
port 88 nsew signal output
flabel metal2 s 12898 21601 12954 22401 0 FreeSans 224 90 0 0 Pin_out[12]
port 89 nsew signal output
flabel metal3 s 19457 6808 20257 6928 0 FreeSans 480 0 0 0 Pin_out[13]
port 90 nsew signal output
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 Pin_out[14]
port 91 nsew signal output
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 Pin_out[15]
port 92 nsew signal output
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 Pin_out[1]
port 93 nsew signal output
flabel metal3 s 19457 9528 20257 9648 0 FreeSans 480 0 0 0 Pin_out[2]
port 94 nsew signal output
flabel metal2 s 5170 21601 5226 22401 0 FreeSans 224 90 0 0 Pin_out[3]
port 95 nsew signal output
flabel metal3 s 19457 21768 20257 21888 0 FreeSans 480 0 0 0 Pin_out[4]
port 96 nsew signal output
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 Pin_out[5]
port 97 nsew signal output
flabel metal2 s 8390 21601 8446 22401 0 FreeSans 224 90 0 0 Pin_out[6]
port 98 nsew signal output
flabel metal3 s 19457 13608 20257 13728 0 FreeSans 480 0 0 0 Pin_out[7]
port 99 nsew signal output
flabel metal3 s 19457 18368 20257 18488 0 FreeSans 480 0 0 0 Pin_out[8]
port 100 nsew signal output
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 Pin_out[9]
port 101 nsew signal output
flabel metal4 s 3004 2128 3324 20176 0 FreeSans 1920 90 0 0 VGND
port 102 nsew ground bidirectional
flabel metal5 s 1056 4076 19184 4396 0 FreeSans 2560 0 0 0 VGND
port 102 nsew ground bidirectional
flabel metal4 s 2344 2128 2664 20176 0 FreeSans 1920 90 0 0 VPWR
port 103 nsew power bidirectional
flabel metal5 s 1056 3416 19184 3736 0 FreeSans 2560 0 0 0 VPWR
port 103 nsew power bidirectional
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 clk
port 104 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 reset
port 105 nsew signal input
rlabel metal1 10120 19584 10120 19584 0 VGND
rlabel metal1 10120 20128 10120 20128 0 VPWR
rlabel metal1 10994 20026 10994 20026 0 Data_in[0]
rlabel metal2 18814 7633 18814 7633 0 Data_in[10]
rlabel metal2 18814 4301 18814 4301 0 Data_in[11]
rlabel metal2 14306 20859 14306 20859 0 Data_in[12]
rlabel metal2 18814 5423 18814 5423 0 Data_in[13]
rlabel metal3 1096 5508 1096 5508 0 Data_in[14]
rlabel metal1 1334 12954 1334 12954 0 Data_in[15]
rlabel metal2 14214 1520 14214 1520 0 Data_in[1]
rlabel metal2 18814 15181 18814 15181 0 Data_in[2]
rlabel metal3 1050 16388 1050 16388 0 Data_in[3]
rlabel metal2 18078 19737 18078 19737 0 Data_in[4]
rlabel metal2 18814 10353 18814 10353 0 Data_in[5]
rlabel metal2 9798 20859 9798 20859 0 Data_in[6]
rlabel metal2 17802 20587 17802 20587 0 Data_in[7]
rlabel metal2 18078 19023 18078 19023 0 Data_in[8]
rlabel metal2 10350 1520 10350 1520 0 Data_in[9]
rlabel metal3 1188 12308 1188 12308 0 Data_out[0]
rlabel metal2 18538 2601 18538 2601 0 Data_out[10]
rlabel metal2 15502 1588 15502 1588 0 Data_out[11]
rlabel metal1 10764 19822 10764 19822 0 Data_out[12]
rlabel metal2 17710 1921 17710 1921 0 Data_out[13]
rlabel metal3 751 2788 751 2788 0 Data_out[14]
rlabel metal3 866 14348 866 14348 0 Data_out[15]
rlabel metal2 10994 1588 10994 1588 0 Data_out[1]
rlabel metal2 18814 11033 18814 11033 0 Data_out[2]
rlabel metal3 751 18428 751 18428 0 Data_out[3]
rlabel metal2 18814 12903 18814 12903 0 Data_out[4]
rlabel metal2 7774 1588 7774 1588 0 Data_out[5]
rlabel metal2 6762 20757 6762 20757 0 Data_out[6]
rlabel metal1 18860 14994 18860 14994 0 Data_out[7]
rlabel metal2 14950 20757 14950 20757 0 Data_out[8]
rlabel metal2 7130 1588 7130 1588 0 Data_out[9]
rlabel metal3 751 4148 751 4148 0 Enable
rlabel metal2 7222 20757 7222 20757 0 Function[0]
rlabel metal2 18262 1241 18262 1241 0 Function[10]
rlabel metal2 17986 1581 17986 1581 0 Function[11]
rlabel metal1 13800 19822 13800 19822 0 Function[12]
rlabel metal2 18814 6239 18814 6239 0 Function[13]
rlabel metal3 1142 4828 1142 4828 0 Function[14]
rlabel metal3 751 15708 751 15708 0 Function[15]
rlabel metal2 12282 1588 12282 1588 0 Function[1]
rlabel metal2 18814 12257 18814 12257 0 Function[2]
rlabel metal3 751 17748 751 17748 0 Function[3]
rlabel metal2 18814 17017 18814 17017 0 Function[4]
rlabel metal3 751 10268 751 10268 0 Function[5]
rlabel metal2 5934 20757 5934 20757 0 Function[6]
rlabel metal2 18814 15895 18814 15895 0 Function[7]
rlabel metal2 16238 20757 16238 20757 0 Function[8]
rlabel metal2 5842 1588 5842 1588 0 Function[9]
rlabel metal1 1380 7514 1380 7514 0 IRQ_INT[0]
rlabel metal3 751 8908 751 8908 0 IRQ_INT[1]
rlabel metal1 1380 8058 1380 8058 0 IRQ_PIN_CHANGE
rlabel metal3 751 9588 751 9588 0 Int_Mask[0]
rlabel metal3 1050 10948 1050 10948 0 Int_Mask[1]
rlabel metal1 9338 18768 9338 18768 0 PIN_DATA[0]
rlabel metal1 17434 5134 17434 5134 0 PIN_DATA[10]
rlabel metal2 17618 4165 17618 4165 0 PIN_DATA[11]
rlabel metal2 12335 21692 12335 21692 0 PIN_DATA[12]
rlabel metal2 17434 8041 17434 8041 0 PIN_DATA[13]
rlabel metal3 1717 6868 1717 6868 0 PIN_DATA[14]
rlabel metal1 4830 13498 4830 13498 0 PIN_DATA[15]
rlabel metal1 12650 4080 12650 4080 0 PIN_DATA[1]
rlabel metal2 17526 11373 17526 11373 0 PIN_DATA[2]
rlabel metal1 2438 17204 2438 17204 0 PIN_DATA[3]
rlabel metal2 17618 17119 17618 17119 0 PIN_DATA[4]
rlabel metal1 9844 7174 9844 7174 0 PIN_DATA[5]
rlabel metal2 7590 19975 7590 19975 0 PIN_DATA[6]
rlabel metal1 17526 14926 17526 14926 0 PIN_DATA[7]
rlabel metal2 16606 17697 16606 17697 0 PIN_DATA[8]
rlabel metal2 8464 2516 8464 2516 0 PIN_DATA[9]
rlabel metal3 751 6188 751 6188 0 Pin_Change_Mask[14]
rlabel metal3 1096 13668 1096 13668 0 Pin_Change_Mask[15]
rlabel metal2 11730 20859 11730 20859 0 Pin_out[0]
rlabel metal2 18538 8857 18538 8857 0 Pin_out[10]
rlabel metal2 18814 3043 18814 3043 0 Pin_out[11]
rlabel metal2 13018 20859 13018 20859 0 Pin_out[12]
rlabel metal3 19190 6868 19190 6868 0 Pin_out[13]
rlabel metal2 6486 1520 6486 1520 0 Pin_out[14]
rlabel metal3 1050 15028 1050 15028 0 Pin_out[15]
rlabel metal2 13570 1520 13570 1520 0 Pin_out[1]
rlabel metal2 18814 9367 18814 9367 0 Pin_out[2]
rlabel metal2 5290 20859 5290 20859 0 Pin_out[3]
rlabel metal2 17526 20927 17526 20927 0 Pin_out[4]
rlabel metal2 11638 1656 11638 1656 0 Pin_out[5]
rlabel metal2 8510 20859 8510 20859 0 Pin_out[6]
rlabel metal2 18814 13855 18814 13855 0 Pin_out[7]
rlabel via2 18814 18411 18814 18411 0 Pin_out[8]
rlabel metal2 9062 1520 9062 1520 0 Pin_out[9]
rlabel metal2 1794 5406 1794 5406 0 _000_
rlabel metal1 3128 7514 3128 7514 0 _001_
rlabel metal2 4002 3230 4002 3230 0 _002_
rlabel metal1 2392 12954 2392 12954 0 _003_
rlabel metal2 4186 10574 4186 10574 0 _004_
rlabel metal2 1702 14688 1702 14688 0 _005_
rlabel metal1 7406 15028 7406 15028 0 _006_
rlabel metal2 16606 6120 16606 6120 0 _007_
rlabel metal2 16974 3060 16974 3060 0 _008_
rlabel metal1 10672 18938 10672 18938 0 _009_
rlabel metal1 16054 7276 16054 7276 0 _010_
rlabel metal1 11132 2890 11132 2890 0 _011_
rlabel metal2 16882 10540 16882 10540 0 _012_
rlabel metal1 2622 18258 2622 18258 0 _013_
rlabel metal2 17342 15198 17342 15198 0 _014_
rlabel metal1 8694 5814 8694 5814 0 _015_
rlabel metal2 6486 18904 6486 18904 0 _016_
rlabel metal1 16238 13362 16238 13362 0 _017_
rlabel metal1 15962 19210 15962 19210 0 _018_
rlabel metal1 6854 2890 6854 2890 0 _019_
rlabel metal1 10817 5270 10817 5270 0 _020_
rlabel metal1 3956 18938 3956 18938 0 _021_
rlabel metal2 4094 16286 4094 16286 0 _022_
rlabel metal1 18032 11322 18032 11322 0 _023_
rlabel metal2 15686 10846 15686 10846 0 _024_
rlabel metal2 17526 15912 17526 15912 0 _025_
rlabel metal2 14582 15946 14582 15946 0 _026_
rlabel metal2 2806 16320 2806 16320 0 _027_
rlabel metal1 3358 18394 3358 18394 0 _028_
rlabel metal2 9614 5032 9614 5032 0 _029_
rlabel metal2 9062 7582 9062 7582 0 _030_
rlabel metal2 18446 16762 18446 16762 0 _031_
rlabel metal1 13340 15674 13340 15674 0 _032_
rlabel metal1 7268 19142 7268 19142 0 _033_
rlabel metal2 6118 16762 6118 16762 0 _034_
rlabel metal1 11415 8874 11415 8874 0 _035_
rlabel metal1 9299 6358 9299 6358 0 _036_
rlabel metal1 18039 13226 18039 13226 0 _037_
rlabel metal2 16054 13906 16054 13906 0 _038_
rlabel metal2 8602 17374 8602 17374 0 _039_
rlabel metal2 5658 18904 5658 18904 0 _040_
rlabel metal2 16974 19176 16974 19176 0 _041_
rlabel metal1 14812 17306 14812 17306 0 _042_
rlabel metal2 18078 14178 18078 14178 0 _043_
rlabel metal1 14260 14246 14260 14246 0 _044_
rlabel metal2 9798 3298 9798 3298 0 _045_
rlabel metal1 8326 2618 8326 2618 0 _046_
rlabel metal1 7084 4998 7084 4998 0 _047_
rlabel metal2 17710 18088 17710 18088 0 _048_
rlabel metal1 15364 18122 15364 18122 0 _049_
rlabel metal1 17388 9146 17388 9146 0 _050_
rlabel metal1 14115 5610 14115 5610 0 _051_
rlabel metal1 9568 18938 9568 18938 0 _052_
rlabel metal1 8011 15402 8011 15402 0 _053_
rlabel metal1 17296 2618 17296 2618 0 _054_
rlabel metal1 15456 4998 15456 4998 0 _055_
rlabel metal1 18078 5338 18078 5338 0 _056_
rlabel metal1 13899 6766 13899 6766 0 _057_
rlabel metal1 11316 18938 11316 18938 0 _058_
rlabel metal1 12427 16490 12427 16490 0 _059_
rlabel metal1 18492 3706 18492 3706 0 _060_
rlabel metal2 15870 3298 15870 3298 0 _061_
rlabel metal1 16836 6426 16836 6426 0 _062_
rlabel metal1 15923 8874 15923 8874 0 _063_
rlabel metal1 13064 18394 13064 18394 0 _064_
rlabel metal1 10994 17510 10994 17510 0 _065_
rlabel metal1 7091 6698 7091 6698 0 _066_
rlabel metal2 13018 12002 13018 12002 0 _067_
rlabel metal1 2300 8058 2300 8058 0 _068_
rlabel metal1 5435 3094 5435 3094 0 _069_
rlabel metal1 5803 5610 5803 5610 0 _070_
rlabel metal2 2898 4998 2898 4998 0 _071_
rlabel metal2 2438 6562 2438 6562 0 _072_
rlabel metal1 5520 7514 5520 7514 0 _073_
rlabel metal1 2944 9146 2944 9146 0 _074_
rlabel metal1 2346 10234 2346 10234 0 _075_
rlabel metal1 7275 11050 7275 11050 0 _076_
rlabel metal1 5619 9622 5619 9622 0 _077_
rlabel metal2 2806 14790 2806 14790 0 _078_
rlabel metal1 6079 13226 6079 13226 0 _079_
rlabel metal2 3174 13464 3174 13464 0 _080_
rlabel metal1 5205 4114 5205 4114 0 _081_
rlabel metal2 2162 11560 2162 11560 0 _082_
rlabel metal1 5205 10710 5205 10710 0 _083_
rlabel metal1 7091 3434 7091 3434 0 _084_
rlabel metal1 10771 15402 10771 15402 0 _085_
rlabel metal1 8556 15674 8556 15674 0 _086_
rlabel metal2 5750 15198 5750 15198 0 _087_
rlabel metal1 12190 2618 12190 2618 0 _088_
rlabel metal2 12558 5406 12558 5406 0 _089_
rlabel metal1 18308 8058 18308 8058 0 _090_
rlabel metal1 14306 7718 14306 7718 0 _091_
rlabel metal1 18315 9962 18315 9962 0 _092_
rlabel metal2 15134 12002 15134 12002 0 _093_
rlabel metal2 13478 3672 13478 3672 0 _094_
rlabel metal1 11132 4794 11132 4794 0 _095_
rlabel metal1 17204 11322 17204 11322 0 _096_
rlabel metal2 15226 10404 15226 10404 0 _097_
rlabel metal1 2024 16626 2024 16626 0 _098_
rlabel metal2 2346 18530 2346 18530 0 _099_
rlabel metal2 17342 16796 17342 16796 0 _100_
rlabel metal2 14122 15572 14122 15572 0 _101_
rlabel metal1 9798 9010 9798 9010 0 _102_
rlabel metal1 8924 5882 8924 5882 0 _103_
rlabel metal1 7912 17238 7912 17238 0 _104_
rlabel metal1 5106 18394 5106 18394 0 _105_
rlabel metal2 17342 14620 17342 14620 0 _106_
rlabel metal2 13202 12954 13202 12954 0 _107_
rlabel metal1 9016 3434 9016 3434 0 _108_
rlabel metal2 16974 18020 16974 18020 0 _109_
rlabel metal2 14674 18530 14674 18530 0 _110_
rlabel metal1 8878 18938 8878 18938 0 _111_
rlabel metal2 7222 15232 7222 15232 0 _112_
rlabel metal1 17112 5338 17112 5338 0 _113_
rlabel metal1 13287 6970 13287 6970 0 _114_
rlabel metal1 17296 3706 17296 3706 0 _115_
rlabel metal2 14398 3672 14398 3672 0 _116_
rlabel metal2 12190 18530 12190 18530 0 _117_
rlabel metal2 9890 17374 9890 17374 0 _118_
rlabel metal1 6111 6970 6111 6970 0 _119_
rlabel metal1 4335 7786 4335 7786 0 _120_
rlabel metal1 6256 10778 6256 10778 0 _121_
rlabel metal1 3726 4046 3726 4046 0 _122_
rlabel metal1 5198 11288 5198 11288 0 _123_
rlabel metal2 5842 3740 5842 3740 0 _124_
rlabel metal1 3956 14586 3956 14586 0 _125_
rlabel metal1 17112 8058 17112 8058 0 _126_
rlabel metal2 14674 7650 14674 7650 0 _127_
rlabel metal2 12282 3808 12282 3808 0 _128_
rlabel metal1 5244 11118 5244 11118 0 _129_
rlabel metal1 2438 5644 2438 5644 0 _130_
rlabel metal1 4324 11050 4324 11050 0 _131_
rlabel metal1 4324 7514 4324 7514 0 _132_
rlabel metal1 4370 8602 4370 8602 0 _133_
rlabel metal2 2346 5780 2346 5780 0 _134_
rlabel metal1 4094 11696 4094 11696 0 _135_
rlabel metal1 11178 17306 11178 17306 0 _136_
rlabel metal1 12696 18261 12696 18261 0 _137_
rlabel metal1 16008 3706 16008 3706 0 _138_
rlabel metal2 17710 3978 17710 3978 0 _139_
rlabel metal2 14490 6528 14490 6528 0 _140_
rlabel metal2 17526 5678 17526 5678 0 _141_
rlabel metal1 7452 15130 7452 15130 0 _142_
rlabel metal2 9430 19210 9430 19210 0 _143_
rlabel metal1 15180 18394 15180 18394 0 _144_
rlabel metal2 16514 18122 16514 18122 0 _145_
rlabel metal2 8326 3740 8326 3740 0 _146_
rlabel metal1 13846 13328 13846 13328 0 _147_
rlabel metal1 17756 14926 17756 14926 0 _148_
rlabel metal1 5888 18394 5888 18394 0 _149_
rlabel metal1 7774 18190 7774 18190 0 _150_
rlabel metal2 9338 6154 9338 6154 0 _151_
rlabel metal1 9292 8602 9292 8602 0 _152_
rlabel metal2 14490 15776 14490 15776 0 _153_
rlabel metal1 17848 17102 17848 17102 0 _154_
rlabel metal1 2806 18394 2806 18394 0 _155_
rlabel metal1 2392 17102 2392 17102 0 _156_
rlabel metal1 15548 10030 15548 10030 0 _157_
rlabel metal2 17618 11594 17618 11594 0 _158_
rlabel metal1 11040 4454 11040 4454 0 _159_
rlabel metal1 12466 4148 12466 4148 0 _160_
rlabel metal1 15134 7514 15134 7514 0 _161_
rlabel metal1 17526 7820 17526 7820 0 _162_
rlabel metal1 4048 14518 4048 14518 0 _163_
rlabel metal1 3910 14314 3910 14314 0 _164_
rlabel metal1 7176 3706 7176 3706 0 _165_
rlabel metal2 4186 11679 4186 11679 0 _166_
rlabel metal1 4876 11186 4876 11186 0 _167_
rlabel metal1 4554 11322 4554 11322 0 _168_
rlabel metal1 5152 11186 5152 11186 0 _169_
rlabel metal1 2254 4046 2254 4046 0 _170_
rlabel metal1 3496 4114 3496 4114 0 _171_
rlabel metal1 4094 6766 4094 6766 0 _172_
rlabel metal2 4186 8160 4186 8160 0 _173_
rlabel metal2 4094 7004 4094 7004 0 _174_
rlabel metal2 4002 7446 4002 7446 0 _175_
rlabel metal2 3542 5508 3542 5508 0 _176_
rlabel metal1 3634 12818 3634 12818 0 _177_
rlabel metal1 5336 5270 5336 5270 0 _178_
rlabel metal1 5520 13974 5520 13974 0 _179_
rlabel metal2 9522 16252 9522 16252 0 _180_
rlabel metal1 12144 4658 12144 4658 0 _181_
rlabel metal1 15916 11730 15916 11730 0 _182_
rlabel metal1 4094 16694 4094 16694 0 _183_
rlabel metal2 16238 15980 16238 15980 0 _184_
rlabel metal1 9614 6902 9614 6902 0 _185_
rlabel metal2 6762 17986 6762 17986 0 _186_
rlabel metal2 15686 13940 15686 13940 0 _187_
rlabel metal1 15640 17306 15640 17306 0 _188_
rlabel metal1 7636 4114 7636 4114 0 _189_
rlabel metal2 15042 5780 15042 5780 0 _190_
rlabel metal2 16422 4454 16422 4454 0 _191_
rlabel metal2 11914 17476 11914 17476 0 _192_
rlabel metal1 15962 8058 15962 8058 0 _193_
rlabel metal3 1395 19108 1395 19108 0 clk
rlabel metal2 12558 7990 12558 7990 0 clknet_0_clk
rlabel metal1 1472 5202 1472 5202 0 clknet_3_0__leaf_clk
rlabel metal1 1702 9554 1702 9554 0 clknet_3_1__leaf_clk
rlabel metal2 17066 3706 17066 3706 0 clknet_3_2__leaf_clk
rlabel metal2 16698 8976 16698 8976 0 clknet_3_3__leaf_clk
rlabel metal1 2714 19380 2714 19380 0 clknet_3_4__leaf_clk
rlabel metal2 1702 17680 1702 17680 0 clknet_3_5__leaf_clk
rlabel metal1 14030 12274 14030 12274 0 clknet_3_6__leaf_clk
rlabel metal2 12650 17782 12650 17782 0 clknet_3_7__leaf_clk
rlabel metal1 1978 5678 1978 5678 0 gpio_instance_14.Data_in
rlabel metal1 4140 5610 4140 5610 0 gpio_instance_14.Function
rlabel metal1 1932 7854 1932 7854 0 gpio_instance_14.IRQ_INT
rlabel metal1 7084 7378 7084 7378 0 gpio_instance_14.PIN_DATA_prev
rlabel metal1 5842 2992 5842 2992 0 gpio_instance_14.Pin_out
rlabel metal1 12466 5712 12466 5712 0 gpio_instance_14.enable_reg
rlabel metal1 5045 5202 5045 5202 0 gpio_instance_14.function_reg
rlabel metal1 3956 9350 3956 9350 0 gpio_instance_14.int_mask_reg\[0\]
rlabel metal2 3910 10948 3910 10948 0 gpio_instance_14.int_mask_reg\[1\]
rlabel metal2 4830 7548 4830 7548 0 gpio_instance_14.irq_detected
rlabel metal1 3358 6188 3358 6188 0 gpio_instance_14.pin_change_mask_reg
rlabel metal1 5336 4250 5336 4250 0 gpio_instance_14.pin_value
rlabel metal1 1840 13294 1840 13294 0 gpio_instance_15.Data_in
rlabel metal2 4646 13532 4646 13532 0 gpio_instance_15.Function
rlabel metal1 1978 8976 1978 8976 0 gpio_instance_15.IRQ_INT
rlabel via1 6854 10982 6854 10982 0 gpio_instance_15.PIN_DATA_prev
rlabel metal1 3312 15130 3312 15130 0 gpio_instance_15.Pin_out
rlabel metal1 6072 13498 6072 13498 0 gpio_instance_15.function_reg
rlabel metal2 5014 11152 5014 11152 0 gpio_instance_15.irq_detected
rlabel metal2 3174 11390 3174 11390 0 gpio_instance_15.pin_change_mask_reg
rlabel via1 5566 14314 5566 14314 0 gpio_instance_15.pin_value
rlabel metal1 9338 19788 9338 19788 0 gpio_pins_0_13\[0\].gpio_instance.Data_in
rlabel metal1 11178 15674 11178 15674 0 gpio_pins_0_13\[0\].gpio_instance.Pin_out
rlabel metal2 9246 16388 9246 16388 0 gpio_pins_0_13\[0\].gpio_instance.function_reg
rlabel metal1 8096 15674 8096 15674 0 gpio_pins_0_13\[0\].gpio_instance.pin_value
rlabel metal1 18354 6290 18354 6290 0 gpio_pins_0_13\[10\].gpio_instance.Data_in
rlabel metal1 18584 9554 18584 9554 0 gpio_pins_0_13\[10\].gpio_instance.Pin_out
rlabel via1 14766 5202 14766 5202 0 gpio_pins_0_13\[10\].gpio_instance.function_reg
rlabel viali 14582 6755 14582 6755 0 gpio_pins_0_13\[10\].gpio_instance.pin_value
rlabel metal2 18814 3740 18814 3740 0 gpio_pins_0_13\[11\].gpio_instance.Data_in
rlabel metal1 18538 2992 18538 2992 0 gpio_pins_0_13\[11\].gpio_instance.Pin_out
rlabel viali 16330 4590 16330 4590 0 gpio_pins_0_13\[11\].gpio_instance.function_reg
rlabel metal2 15870 3876 15870 3876 0 gpio_pins_0_13\[11\].gpio_instance.pin_value
rlabel metal2 13662 19142 13662 19142 0 gpio_pins_0_13\[12\].gpio_instance.Data_in
rlabel metal1 13110 19380 13110 19380 0 gpio_pins_0_13\[12\].gpio_instance.Pin_out
rlabel metal2 12466 16762 12466 16762 0 gpio_pins_0_13\[12\].gpio_instance.function_reg
rlabel metal1 10902 17680 10902 17680 0 gpio_pins_0_13\[12\].gpio_instance.pin_value
rlabel metal2 18170 8058 18170 8058 0 gpio_pins_0_13\[13\].gpio_instance.Data_in
rlabel metal1 18170 6800 18170 6800 0 gpio_pins_0_13\[13\].gpio_instance.Pin_out
rlabel via1 16054 7854 16054 7854 0 gpio_pins_0_13\[13\].gpio_instance.function_reg
rlabel metal1 15824 7718 15824 7718 0 gpio_pins_0_13\[13\].gpio_instance.pin_value
rlabel metal2 13754 3196 13754 3196 0 gpio_pins_0_13\[1\].gpio_instance.Data_in
rlabel metal1 13340 3026 13340 3026 0 gpio_pins_0_13\[1\].gpio_instance.Pin_out
rlabel metal2 13294 5474 13294 5474 0 gpio_pins_0_13\[1\].gpio_instance.function_reg
rlabel metal2 10718 4794 10718 4794 0 gpio_pins_0_13\[1\].gpio_instance.pin_value
rlabel metal1 18446 12206 18446 12206 0 gpio_pins_0_13\[2\].gpio_instance.Data_in
rlabel metal2 18354 10438 18354 10438 0 gpio_pins_0_13\[2\].gpio_instance.Pin_out
rlabel metal1 15625 11730 15625 11730 0 gpio_pins_0_13\[2\].gpio_instance.function_reg
rlabel metal1 15962 10778 15962 10778 0 gpio_pins_0_13\[2\].gpio_instance.pin_value
rlabel metal1 2070 16116 2070 16116 0 gpio_pins_0_13\[3\].gpio_instance.Data_in
rlabel metal1 4600 19346 4600 19346 0 gpio_pins_0_13\[3\].gpio_instance.Pin_out
rlabel metal2 4922 16354 4922 16354 0 gpio_pins_0_13\[3\].gpio_instance.function_reg
rlabel metal2 3542 17884 3542 17884 0 gpio_pins_0_13\[3\].gpio_instance.pin_value
rlabel metal1 18354 17204 18354 17204 0 gpio_pins_0_13\[4\].gpio_instance.Data_in
rlabel metal1 18492 16218 18492 16218 0 gpio_pins_0_13\[4\].gpio_instance.Pin_out
rlabel metal1 14628 15674 14628 15674 0 gpio_pins_0_13\[4\].gpio_instance.function_reg
rlabel metal1 14490 14994 14490 14994 0 gpio_pins_0_13\[4\].gpio_instance.pin_value
rlabel metal1 10626 8806 10626 8806 0 gpio_pins_0_13\[5\].gpio_instance.Data_in
rlabel metal1 11220 3026 11220 3026 0 gpio_pins_0_13\[5\].gpio_instance.Pin_out
rlabel metal1 9369 6766 9369 6766 0 gpio_pins_0_13\[5\].gpio_instance.function_reg
rlabel metal1 9476 6426 9476 6426 0 gpio_pins_0_13\[5\].gpio_instance.pin_value
rlabel metal2 9246 17782 9246 17782 0 gpio_pins_0_13\[6\].gpio_instance.Data_in
rlabel metal1 8004 18734 8004 18734 0 gpio_pins_0_13\[6\].gpio_instance.Pin_out
rlabel metal2 6486 17204 6486 17204 0 gpio_pins_0_13\[6\].gpio_instance.function_reg
rlabel metal2 6026 18428 6026 18428 0 gpio_pins_0_13\[6\].gpio_instance.pin_value
rlabel metal2 18262 17408 18262 17408 0 gpio_pins_0_13\[7\].gpio_instance.Data_in
rlabel metal1 18446 13328 18446 13328 0 gpio_pins_0_13\[7\].gpio_instance.Pin_out
rlabel metal1 15993 12818 15993 12818 0 gpio_pins_0_13\[7\].gpio_instance.function_reg
rlabel metal1 15088 12954 15088 12954 0 gpio_pins_0_13\[7\].gpio_instance.pin_value
rlabel metal1 18308 18734 18308 18734 0 gpio_pins_0_13\[8\].gpio_instance.Data_in
rlabel metal2 18446 18938 18446 18938 0 gpio_pins_0_13\[8\].gpio_instance.Pin_out
rlabel via1 15226 17170 15226 17170 0 gpio_pins_0_13\[8\].gpio_instance.function_reg
rlabel metal1 15640 18258 15640 18258 0 gpio_pins_0_13\[8\].gpio_instance.pin_value
rlabel metal2 10718 3910 10718 3910 0 gpio_pins_0_13\[9\].gpio_instance.Data_in
rlabel metal1 8970 2992 8970 2992 0 gpio_pins_0_13\[9\].gpio_instance.Pin_out
rlabel metal1 7728 4794 7728 4794 0 gpio_pins_0_13\[9\].gpio_instance.function_reg
rlabel metal1 7268 4046 7268 4046 0 gpio_pins_0_13\[9\].gpio_instance.pin_value
rlabel metal2 7038 13838 7038 13838 0 net1
rlabel metal2 1794 18496 1794 18496 0 net10
rlabel metal1 18584 12954 18584 12954 0 net11
rlabel metal1 8326 2550 8326 2550 0 net12
rlabel metal2 6578 19584 6578 19584 0 net13
rlabel metal1 17250 14042 17250 14042 0 net14
rlabel metal2 14950 19584 14950 19584 0 net15
rlabel metal1 7130 2618 7130 2618 0 net16
rlabel metal2 2070 4318 2070 4318 0 net17
rlabel metal1 7084 16082 7084 16082 0 net18
rlabel metal1 17250 5202 17250 5202 0 net19
rlabel metal2 16514 4046 16514 4046 0 net2
rlabel metal1 17526 3536 17526 3536 0 net20
rlabel via1 12925 19346 12925 19346 0 net21
rlabel metal1 18354 6426 18354 6426 0 net22
rlabel metal2 1978 5372 1978 5372 0 net23
rlabel metal2 1794 15130 1794 15130 0 net24
rlabel metal2 12466 2618 12466 2618 0 net25
rlabel viali 18077 12206 18077 12206 0 net26
rlabel metal1 2208 18054 2208 18054 0 net27
rlabel via1 18185 17170 18185 17170 0 net28
rlabel metal1 9338 8976 9338 8976 0 net29
rlabel metal1 15548 2618 15548 2618 0 net3
rlabel metal2 5750 17986 5750 17986 0 net30
rlabel via1 18169 14994 18169 14994 0 net31
rlabel metal1 16529 18734 16529 18734 0 net32
rlabel metal1 6486 2618 6486 2618 0 net33
rlabel metal1 1886 9622 1886 9622 0 net34
rlabel metal1 1656 10710 1656 10710 0 net35
rlabel metal1 2208 5678 2208 5678 0 net36
rlabel metal1 1748 13770 1748 13770 0 net37
rlabel metal1 2346 4590 2346 4590 0 net38
rlabel metal1 11270 19856 11270 19856 0 net39
rlabel metal2 10534 19176 10534 19176 0 net4
rlabel metal2 18630 7412 18630 7412 0 net40
rlabel metal2 18354 4148 18354 4148 0 net41
rlabel metal1 14168 19482 14168 19482 0 net42
rlabel metal1 18584 5202 18584 5202 0 net43
rlabel metal1 1656 5678 1656 5678 0 net44
rlabel metal2 1610 12988 1610 12988 0 net45
rlabel metal2 14490 2618 14490 2618 0 net46
rlabel metal2 18354 14212 18354 14212 0 net47
rlabel metal1 1518 16762 1518 16762 0 net48
rlabel metal1 18216 19482 18216 19482 0 net49
rlabel metal1 17480 2618 17480 2618 0 net5
rlabel metal2 17986 9962 17986 9962 0 net50
rlabel metal1 9706 18394 9706 18394 0 net51
rlabel metal1 17618 19788 17618 19788 0 net52
rlabel metal1 18032 18734 18032 18734 0 net53
rlabel metal1 10442 2822 10442 2822 0 net54
rlabel metal1 2070 7378 2070 7378 0 net55
rlabel metal1 1702 8942 1702 8942 0 net56
rlabel metal1 1656 7854 1656 7854 0 net57
rlabel metal2 11730 19652 11730 19652 0 net58
rlabel metal2 18354 9146 18354 9146 0 net59
rlabel metal1 1656 3162 1656 3162 0 net6
rlabel metal2 18630 2618 18630 2618 0 net60
rlabel metal2 13294 19652 13294 19652 0 net61
rlabel metal2 18354 7174 18354 7174 0 net62
rlabel metal1 6394 2822 6394 2822 0 net63
rlabel metal1 1978 15470 1978 15470 0 net64
rlabel metal2 13846 2618 13846 2618 0 net65
rlabel metal2 18630 9690 18630 9690 0 net66
rlabel metal2 4922 19652 4922 19652 0 net67
rlabel metal1 17342 19856 17342 19856 0 net68
rlabel metal1 11776 2822 11776 2822 0 net69
rlabel metal1 1748 14042 1748 14042 0 net7
rlabel metal1 8464 18938 8464 18938 0 net70
rlabel metal2 18630 13702 18630 13702 0 net71
rlabel metal2 18630 18428 18630 18428 0 net72
rlabel metal1 9246 2822 9246 2822 0 net73
rlabel metal2 11040 3094 11040 3094 0 net8
rlabel metal1 17618 11050 17618 11050 0 net9
rlabel metal3 751 3468 751 3468 0 reset
<< properties >>
string FIXED_BBOX 0 0 20257 22401
<< end >>
