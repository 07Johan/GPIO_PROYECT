module gpio_vector (Enable,
    IRQ_PIN_CHANGE,
    clk,
    reset,
    Data_in,
    Data_out,
    Function,
    IRQ_INT,
    Int_Mask,
    PIN_DATA,
    Pin_Change_Mask,
    Pin_out);
 input Enable;
 output IRQ_PIN_CHANGE;
 input clk;
 input reset;
 output [15:0] Data_in;
 input [15:0] Data_out;
 input [15:0] Function;
 output [1:0] IRQ_INT;
 input [1:0] Int_Mask;
 inout [15:0] PIN_DATA;
 input [15:0] Pin_Change_Mask;
 output [15:0] Pin_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire \gpio_instance_14.Data_in ;
 wire \gpio_instance_14.Function ;
 wire \gpio_instance_14.IRQ_INT ;
 wire \gpio_instance_14.PIN_DATA_prev ;
 wire \gpio_instance_14.Pin_out ;
 wire \gpio_instance_14.enable_reg ;
 wire \gpio_instance_14.function_reg ;
 wire \gpio_instance_14.int_mask_reg[0] ;
 wire \gpio_instance_14.int_mask_reg[1] ;
 wire \gpio_instance_14.irq_detected ;
 wire \gpio_instance_14.pin_change_mask_reg ;
 wire \gpio_instance_14.pin_value ;
 wire \gpio_instance_15.Data_in ;
 wire \gpio_instance_15.Function ;
 wire \gpio_instance_15.IRQ_INT ;
 wire \gpio_instance_15.PIN_DATA_prev ;
 wire \gpio_instance_15.Pin_out ;
 wire \gpio_instance_15.function_reg ;
 wire \gpio_instance_15.irq_detected ;
 wire \gpio_instance_15.pin_change_mask_reg ;
 wire \gpio_instance_15.pin_value ;
 wire \gpio_pins_0_13[0].gpio_instance.Data_in ;
 wire \gpio_pins_0_13[0].gpio_instance.Pin_out ;
 wire \gpio_pins_0_13[0].gpio_instance.function_reg ;
 wire \gpio_pins_0_13[0].gpio_instance.pin_value ;
 wire \gpio_pins_0_13[10].gpio_instance.Data_in ;
 wire \gpio_pins_0_13[10].gpio_instance.Pin_out ;
 wire \gpio_pins_0_13[10].gpio_instance.function_reg ;
 wire \gpio_pins_0_13[10].gpio_instance.pin_value ;
 wire \gpio_pins_0_13[11].gpio_instance.Data_in ;
 wire \gpio_pins_0_13[11].gpio_instance.Pin_out ;
 wire \gpio_pins_0_13[11].gpio_instance.function_reg ;
 wire \gpio_pins_0_13[11].gpio_instance.pin_value ;
 wire \gpio_pins_0_13[12].gpio_instance.Data_in ;
 wire \gpio_pins_0_13[12].gpio_instance.Pin_out ;
 wire \gpio_pins_0_13[12].gpio_instance.function_reg ;
 wire \gpio_pins_0_13[12].gpio_instance.pin_value ;
 wire \gpio_pins_0_13[13].gpio_instance.Data_in ;
 wire \gpio_pins_0_13[13].gpio_instance.Pin_out ;
 wire \gpio_pins_0_13[13].gpio_instance.function_reg ;
 wire \gpio_pins_0_13[13].gpio_instance.pin_value ;
 wire \gpio_pins_0_13[1].gpio_instance.Data_in ;
 wire \gpio_pins_0_13[1].gpio_instance.Pin_out ;
 wire \gpio_pins_0_13[1].gpio_instance.function_reg ;
 wire \gpio_pins_0_13[1].gpio_instance.pin_value ;
 wire \gpio_pins_0_13[2].gpio_instance.Data_in ;
 wire \gpio_pins_0_13[2].gpio_instance.Pin_out ;
 wire \gpio_pins_0_13[2].gpio_instance.function_reg ;
 wire \gpio_pins_0_13[2].gpio_instance.pin_value ;
 wire \gpio_pins_0_13[3].gpio_instance.Data_in ;
 wire \gpio_pins_0_13[3].gpio_instance.Pin_out ;
 wire \gpio_pins_0_13[3].gpio_instance.function_reg ;
 wire \gpio_pins_0_13[3].gpio_instance.pin_value ;
 wire \gpio_pins_0_13[4].gpio_instance.Data_in ;
 wire \gpio_pins_0_13[4].gpio_instance.Pin_out ;
 wire \gpio_pins_0_13[4].gpio_instance.function_reg ;
 wire \gpio_pins_0_13[4].gpio_instance.pin_value ;
 wire \gpio_pins_0_13[5].gpio_instance.Data_in ;
 wire \gpio_pins_0_13[5].gpio_instance.Pin_out ;
 wire \gpio_pins_0_13[5].gpio_instance.function_reg ;
 wire \gpio_pins_0_13[5].gpio_instance.pin_value ;
 wire \gpio_pins_0_13[6].gpio_instance.Data_in ;
 wire \gpio_pins_0_13[6].gpio_instance.Pin_out ;
 wire \gpio_pins_0_13[6].gpio_instance.function_reg ;
 wire \gpio_pins_0_13[6].gpio_instance.pin_value ;
 wire \gpio_pins_0_13[7].gpio_instance.Data_in ;
 wire \gpio_pins_0_13[7].gpio_instance.Pin_out ;
 wire \gpio_pins_0_13[7].gpio_instance.function_reg ;
 wire \gpio_pins_0_13[7].gpio_instance.pin_value ;
 wire \gpio_pins_0_13[8].gpio_instance.Data_in ;
 wire \gpio_pins_0_13[8].gpio_instance.Pin_out ;
 wire \gpio_pins_0_13[8].gpio_instance.function_reg ;
 wire \gpio_pins_0_13[8].gpio_instance.pin_value ;
 wire \gpio_pins_0_13[9].gpio_instance.Data_in ;
 wire \gpio_pins_0_13[9].gpio_instance.Pin_out ;
 wire \gpio_pins_0_13[9].gpio_instance.function_reg ;
 wire \gpio_pins_0_13[9].gpio_instance.pin_value ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sky130_fd_sc_hd__inv_2 _194_ (.A(\gpio_instance_15.irq_detected ),
    .Y(_129_));
 sky130_fd_sc_hd__inv_8 _195_ (.A(net17),
    .Y(_130_));
 sky130_fd_sc_hd__inv_2 _196_ (.A(\gpio_instance_15.PIN_DATA_prev ),
    .Y(_131_));
 sky130_fd_sc_hd__inv_2 _197_ (.A(\gpio_instance_14.irq_detected ),
    .Y(_132_));
 sky130_fd_sc_hd__inv_2 _198_ (.A(\gpio_instance_14.PIN_DATA_prev ),
    .Y(_133_));
 sky130_fd_sc_hd__inv_2 _199_ (.A(net23),
    .Y(_134_));
 sky130_fd_sc_hd__inv_2 _200_ (.A(net24),
    .Y(_135_));
 sky130_fd_sc_hd__inv_2 _201_ (.A(net38),
    .Y(_066_));
 sky130_fd_sc_hd__nand2_1 _202_ (.A(_130_),
    .B(net21),
    .Y(_136_));
 sky130_fd_sc_hd__and3b_1 _203_ (.A_N(net17),
    .B(net21),
    .C(net4),
    .X(_009_));
 sky130_fd_sc_hd__a21o_1 _204_ (.A1(_136_),
    .A2(\gpio_pins_0_13[12].gpio_instance.pin_value ),
    .B1(_009_),
    .X(_118_));
 sky130_fd_sc_hd__nand2b_1 _205_ (.A_N(\gpio_pins_0_13[12].gpio_instance.Data_in ),
    .B(net21),
    .Y(_137_));
 sky130_fd_sc_hd__o211a_1 _206_ (.A1(net21),
    .A2(PIN_DATA[12]),
    .B1(_137_),
    .C1(_130_),
    .X(_117_));
 sky130_fd_sc_hd__nand2_1 _207_ (.A(_130_),
    .B(net20),
    .Y(_138_));
 sky130_fd_sc_hd__and3b_1 _208_ (.A_N(net17),
    .B(net20),
    .C(net3),
    .X(_008_));
 sky130_fd_sc_hd__a21o_1 _209_ (.A1(_138_),
    .A2(\gpio_pins_0_13[11].gpio_instance.pin_value ),
    .B1(_008_),
    .X(_116_));
 sky130_fd_sc_hd__nand2b_1 _210_ (.A_N(\gpio_pins_0_13[11].gpio_instance.Data_in ),
    .B(net20),
    .Y(_139_));
 sky130_fd_sc_hd__o211a_1 _211_ (.A1(net20),
    .A2(PIN_DATA[11]),
    .B1(_139_),
    .C1(_130_),
    .X(_115_));
 sky130_fd_sc_hd__nand2_1 _212_ (.A(_130_),
    .B(net19),
    .Y(_140_));
 sky130_fd_sc_hd__and3b_1 _213_ (.A_N(net17),
    .B(net19),
    .C(net2),
    .X(_007_));
 sky130_fd_sc_hd__a21o_1 _214_ (.A1(_140_),
    .A2(\gpio_pins_0_13[10].gpio_instance.pin_value ),
    .B1(_007_),
    .X(_114_));
 sky130_fd_sc_hd__nand2b_1 _215_ (.A_N(\gpio_pins_0_13[10].gpio_instance.Data_in ),
    .B(net19),
    .Y(_141_));
 sky130_fd_sc_hd__o211a_1 _216_ (.A1(net19),
    .A2(PIN_DATA[10]),
    .B1(_141_),
    .C1(_130_),
    .X(_113_));
 sky130_fd_sc_hd__nand2_1 _217_ (.A(_130_),
    .B(net18),
    .Y(_142_));
 sky130_fd_sc_hd__and3b_1 _218_ (.A_N(net17),
    .B(net18),
    .C(net1),
    .X(_006_));
 sky130_fd_sc_hd__a21o_1 _219_ (.A1(_142_),
    .A2(\gpio_pins_0_13[0].gpio_instance.pin_value ),
    .B1(_006_),
    .X(_112_));
 sky130_fd_sc_hd__nand2b_1 _220_ (.A_N(\gpio_pins_0_13[0].gpio_instance.Data_in ),
    .B(net18),
    .Y(_143_));
 sky130_fd_sc_hd__o211a_1 _221_ (.A1(net18),
    .A2(PIN_DATA[0]),
    .B1(_143_),
    .C1(_130_),
    .X(_111_));
 sky130_fd_sc_hd__nand2_1 _222_ (.A(_130_),
    .B(net32),
    .Y(_144_));
 sky130_fd_sc_hd__and3b_1 _223_ (.A_N(net17),
    .B(net32),
    .C(net15),
    .X(_018_));
 sky130_fd_sc_hd__a21o_1 _224_ (.A1(_144_),
    .A2(\gpio_pins_0_13[8].gpio_instance.pin_value ),
    .B1(_018_),
    .X(_110_));
 sky130_fd_sc_hd__nand2b_1 _225_ (.A_N(\gpio_pins_0_13[8].gpio_instance.Data_in ),
    .B(net32),
    .Y(_145_));
 sky130_fd_sc_hd__o211a_1 _226_ (.A1(net32),
    .A2(PIN_DATA[8]),
    .B1(_145_),
    .C1(_130_),
    .X(_109_));
 sky130_fd_sc_hd__nand2b_1 _227_ (.A_N(\gpio_pins_0_13[9].gpio_instance.Data_in ),
    .B(net33),
    .Y(_146_));
 sky130_fd_sc_hd__o211a_1 _228_ (.A1(net33),
    .A2(PIN_DATA[9]),
    .B1(_146_),
    .C1(_130_),
    .X(_108_));
 sky130_fd_sc_hd__nand2_1 _229_ (.A(_130_),
    .B(net31),
    .Y(_147_));
 sky130_fd_sc_hd__and3b_1 _230_ (.A_N(net17),
    .B(net31),
    .C(net14),
    .X(_017_));
 sky130_fd_sc_hd__a21o_1 _231_ (.A1(_147_),
    .A2(\gpio_pins_0_13[7].gpio_instance.pin_value ),
    .B1(_017_),
    .X(_107_));
 sky130_fd_sc_hd__nand2b_1 _232_ (.A_N(\gpio_pins_0_13[7].gpio_instance.Data_in ),
    .B(net31),
    .Y(_148_));
 sky130_fd_sc_hd__o211a_1 _233_ (.A1(net31),
    .A2(PIN_DATA[7]),
    .B1(_148_),
    .C1(_130_),
    .X(_106_));
 sky130_fd_sc_hd__nand2_1 _234_ (.A(_130_),
    .B(net30),
    .Y(_149_));
 sky130_fd_sc_hd__and3b_1 _235_ (.A_N(net17),
    .B(net30),
    .C(net13),
    .X(_016_));
 sky130_fd_sc_hd__a21o_1 _236_ (.A1(_149_),
    .A2(\gpio_pins_0_13[6].gpio_instance.pin_value ),
    .B1(_016_),
    .X(_105_));
 sky130_fd_sc_hd__nand2b_1 _237_ (.A_N(\gpio_pins_0_13[6].gpio_instance.Data_in ),
    .B(net30),
    .Y(_150_));
 sky130_fd_sc_hd__o211a_1 _238_ (.A1(net30),
    .A2(PIN_DATA[6]),
    .B1(_150_),
    .C1(_130_),
    .X(_104_));
 sky130_fd_sc_hd__nand2_1 _239_ (.A(_130_),
    .B(net29),
    .Y(_151_));
 sky130_fd_sc_hd__and3b_1 _240_ (.A_N(net17),
    .B(net29),
    .C(net12),
    .X(_015_));
 sky130_fd_sc_hd__a21o_1 _241_ (.A1(_151_),
    .A2(\gpio_pins_0_13[5].gpio_instance.pin_value ),
    .B1(_015_),
    .X(_103_));
 sky130_fd_sc_hd__nand2b_1 _242_ (.A_N(\gpio_pins_0_13[5].gpio_instance.Data_in ),
    .B(net29),
    .Y(_152_));
 sky130_fd_sc_hd__o211a_1 _243_ (.A1(net29),
    .A2(PIN_DATA[5]),
    .B1(_152_),
    .C1(_130_),
    .X(_102_));
 sky130_fd_sc_hd__nand2_1 _244_ (.A(_130_),
    .B(net28),
    .Y(_153_));
 sky130_fd_sc_hd__and3b_1 _245_ (.A_N(net17),
    .B(net28),
    .C(net11),
    .X(_014_));
 sky130_fd_sc_hd__a21o_1 _246_ (.A1(_153_),
    .A2(\gpio_pins_0_13[4].gpio_instance.pin_value ),
    .B1(_014_),
    .X(_101_));
 sky130_fd_sc_hd__nand2b_1 _247_ (.A_N(\gpio_pins_0_13[4].gpio_instance.Data_in ),
    .B(net28),
    .Y(_154_));
 sky130_fd_sc_hd__o211a_1 _248_ (.A1(net28),
    .A2(PIN_DATA[4]),
    .B1(_154_),
    .C1(_130_),
    .X(_100_));
 sky130_fd_sc_hd__nand2_1 _249_ (.A(_130_),
    .B(net27),
    .Y(_155_));
 sky130_fd_sc_hd__and3b_1 _250_ (.A_N(net17),
    .B(net27),
    .C(net10),
    .X(_013_));
 sky130_fd_sc_hd__a21o_1 _251_ (.A1(_155_),
    .A2(\gpio_pins_0_13[3].gpio_instance.pin_value ),
    .B1(_013_),
    .X(_099_));
 sky130_fd_sc_hd__nand2b_1 _252_ (.A_N(\gpio_pins_0_13[3].gpio_instance.Data_in ),
    .B(net27),
    .Y(_156_));
 sky130_fd_sc_hd__o211a_1 _253_ (.A1(net27),
    .A2(PIN_DATA[3]),
    .B1(_156_),
    .C1(_130_),
    .X(_098_));
 sky130_fd_sc_hd__nand2_1 _254_ (.A(_130_),
    .B(net26),
    .Y(_157_));
 sky130_fd_sc_hd__and3b_1 _255_ (.A_N(net17),
    .B(net26),
    .C(net9),
    .X(_012_));
 sky130_fd_sc_hd__a21o_1 _256_ (.A1(_157_),
    .A2(\gpio_pins_0_13[2].gpio_instance.pin_value ),
    .B1(_012_),
    .X(_097_));
 sky130_fd_sc_hd__nand2b_1 _257_ (.A_N(\gpio_pins_0_13[2].gpio_instance.Data_in ),
    .B(net26),
    .Y(_158_));
 sky130_fd_sc_hd__o211a_1 _258_ (.A1(net26),
    .A2(PIN_DATA[2]),
    .B1(_158_),
    .C1(_130_),
    .X(_096_));
 sky130_fd_sc_hd__nand2_1 _259_ (.A(_130_),
    .B(net25),
    .Y(_159_));
 sky130_fd_sc_hd__and3b_1 _260_ (.A_N(net17),
    .B(net25),
    .C(net8),
    .X(_011_));
 sky130_fd_sc_hd__a21o_1 _261_ (.A1(_159_),
    .A2(\gpio_pins_0_13[1].gpio_instance.pin_value ),
    .B1(_011_),
    .X(_095_));
 sky130_fd_sc_hd__nand2b_1 _262_ (.A_N(\gpio_pins_0_13[1].gpio_instance.Data_in ),
    .B(net25),
    .Y(_160_));
 sky130_fd_sc_hd__o211a_1 _263_ (.A1(net25),
    .A2(PIN_DATA[1]),
    .B1(_160_),
    .C1(_130_),
    .X(_128_));
 sky130_fd_sc_hd__nand2_1 _264_ (.A(_130_),
    .B(net22),
    .Y(_161_));
 sky130_fd_sc_hd__and3b_1 _265_ (.A_N(net17),
    .B(net22),
    .C(net5),
    .X(_010_));
 sky130_fd_sc_hd__a21o_1 _266_ (.A1(_161_),
    .A2(\gpio_pins_0_13[13].gpio_instance.pin_value ),
    .B1(_010_),
    .X(_127_));
 sky130_fd_sc_hd__nand2b_1 _267_ (.A_N(\gpio_pins_0_13[13].gpio_instance.Data_in ),
    .B(net22),
    .Y(_162_));
 sky130_fd_sc_hd__o211a_1 _268_ (.A1(net22),
    .A2(PIN_DATA[13]),
    .B1(_162_),
    .C1(_130_),
    .X(_126_));
 sky130_fd_sc_hd__nor2_1 _269_ (.A(net37),
    .B(_135_),
    .Y(\gpio_instance_15.Function ));
 sky130_fd_sc_hd__nor2_1 _270_ (.A(net17),
    .B(net37),
    .Y(_163_));
 sky130_fd_sc_hd__nand2_1 _271_ (.A(net24),
    .B(_163_),
    .Y(_164_));
 sky130_fd_sc_hd__and4bb_1 _272_ (.A_N(net17),
    .B_N(net37),
    .C(net24),
    .D(net7),
    .X(_005_));
 sky130_fd_sc_hd__a21o_1 _273_ (.A1(_164_),
    .A2(\gpio_instance_15.pin_value ),
    .B1(_005_),
    .X(_125_));
 sky130_fd_sc_hd__nand2_1 _274_ (.A(_130_),
    .B(net33),
    .Y(_165_));
 sky130_fd_sc_hd__and3b_1 _275_ (.A_N(net17),
    .B(net33),
    .C(net16),
    .X(_019_));
 sky130_fd_sc_hd__a21o_1 _276_ (.A1(_165_),
    .A2(\gpio_pins_0_13[9].gpio_instance.pin_value ),
    .B1(_019_),
    .X(_124_));
 sky130_fd_sc_hd__and2b_1 _277_ (.A_N(net17),
    .B(\gpio_instance_15.pin_change_mask_reg ),
    .X(_166_));
 sky130_fd_sc_hd__a21boi_1 _278_ (.A1(_131_),
    .A2(\gpio_instance_14.int_mask_reg[0] ),
    .B1_N(PIN_DATA[15]),
    .Y(_167_));
 sky130_fd_sc_hd__a21o_1 _279_ (.A1(\gpio_instance_15.PIN_DATA_prev ),
    .A2(\gpio_instance_14.int_mask_reg[1] ),
    .B1(PIN_DATA[15]),
    .X(_168_));
 sky130_fd_sc_hd__o211ai_1 _280_ (.A1(net37),
    .A2(_135_),
    .B1(_168_),
    .C1(_166_),
    .Y(_169_));
 sky130_fd_sc_hd__o22ai_1 _281_ (.A1(_129_),
    .A2(_130_),
    .B1(_167_),
    .B2(_169_),
    .Y(_123_));
 sky130_fd_sc_hd__nor2_1 _282_ (.A(net36),
    .B(_134_),
    .Y(\gpio_instance_14.Function ));
 sky130_fd_sc_hd__or4bb_1 _283_ (.A(net17),
    .B(net36),
    .C_N(net23),
    .D_N(net6),
    .X(_170_));
 sky130_fd_sc_hd__inv_2 _284_ (.A(_170_),
    .Y(_002_));
 sky130_fd_sc_hd__o31ai_1 _285_ (.A1(net17),
    .A2(net36),
    .A3(_134_),
    .B1(\gpio_instance_14.pin_value ),
    .Y(_171_));
 sky130_fd_sc_hd__nand2_1 _286_ (.A(_170_),
    .B(_171_),
    .Y(_122_));
 sky130_fd_sc_hd__mux2_1 _287_ (.A0(PIN_DATA[15]),
    .A1(\gpio_instance_15.PIN_DATA_prev ),
    .S(net17),
    .X(_121_));
 sky130_fd_sc_hd__and2b_1 _288_ (.A_N(net17),
    .B(\gpio_instance_14.pin_change_mask_reg ),
    .X(_172_));
 sky130_fd_sc_hd__a21boi_1 _289_ (.A1(_133_),
    .A2(\gpio_instance_14.int_mask_reg[0] ),
    .B1_N(PIN_DATA[14]),
    .Y(_173_));
 sky130_fd_sc_hd__a21o_1 _290_ (.A1(\gpio_instance_14.PIN_DATA_prev ),
    .A2(\gpio_instance_14.int_mask_reg[1] ),
    .B1(PIN_DATA[14]),
    .X(_174_));
 sky130_fd_sc_hd__o211ai_1 _291_ (.A1(net36),
    .A2(_134_),
    .B1(_174_),
    .C1(_172_),
    .Y(_175_));
 sky130_fd_sc_hd__o22ai_1 _292_ (.A1(_130_),
    .A2(_132_),
    .B1(_173_),
    .B2(_175_),
    .Y(_120_));
 sky130_fd_sc_hd__mux2_1 _293_ (.A0(PIN_DATA[14]),
    .A1(\gpio_instance_14.PIN_DATA_prev ),
    .S(net17),
    .X(_119_));
 sky130_fd_sc_hd__nand2b_1 _294_ (.A_N(\gpio_instance_14.enable_reg ),
    .B(\gpio_pins_0_13[13].gpio_instance.function_reg ),
    .Y(_193_));
 sky130_fd_sc_hd__nand2b_1 _295_ (.A_N(\gpio_instance_14.enable_reg ),
    .B(\gpio_pins_0_13[12].gpio_instance.function_reg ),
    .Y(_192_));
 sky130_fd_sc_hd__nand2b_1 _296_ (.A_N(\gpio_instance_14.enable_reg ),
    .B(\gpio_pins_0_13[11].gpio_instance.function_reg ),
    .Y(_191_));
 sky130_fd_sc_hd__nand2b_1 _297_ (.A_N(\gpio_instance_14.enable_reg ),
    .B(\gpio_pins_0_13[10].gpio_instance.function_reg ),
    .Y(_190_));
 sky130_fd_sc_hd__nand2b_1 _298_ (.A_N(\gpio_instance_14.enable_reg ),
    .B(\gpio_pins_0_13[9].gpio_instance.function_reg ),
    .Y(_189_));
 sky130_fd_sc_hd__nand2b_1 _299_ (.A_N(\gpio_instance_14.enable_reg ),
    .B(\gpio_pins_0_13[8].gpio_instance.function_reg ),
    .Y(_188_));
 sky130_fd_sc_hd__nand2b_1 _300_ (.A_N(\gpio_instance_14.enable_reg ),
    .B(\gpio_pins_0_13[7].gpio_instance.function_reg ),
    .Y(_187_));
 sky130_fd_sc_hd__nand2b_1 _301_ (.A_N(\gpio_instance_14.enable_reg ),
    .B(\gpio_pins_0_13[6].gpio_instance.function_reg ),
    .Y(_186_));
 sky130_fd_sc_hd__nand2b_1 _302_ (.A_N(\gpio_instance_14.enable_reg ),
    .B(\gpio_pins_0_13[5].gpio_instance.function_reg ),
    .Y(_185_));
 sky130_fd_sc_hd__nand2b_1 _303_ (.A_N(\gpio_instance_14.enable_reg ),
    .B(\gpio_pins_0_13[4].gpio_instance.function_reg ),
    .Y(_184_));
 sky130_fd_sc_hd__nand2b_1 _304_ (.A_N(\gpio_instance_14.enable_reg ),
    .B(\gpio_pins_0_13[3].gpio_instance.function_reg ),
    .Y(_183_));
 sky130_fd_sc_hd__nand2b_1 _305_ (.A_N(\gpio_instance_14.enable_reg ),
    .B(\gpio_pins_0_13[2].gpio_instance.function_reg ),
    .Y(_182_));
 sky130_fd_sc_hd__nand2b_1 _306_ (.A_N(\gpio_instance_14.enable_reg ),
    .B(\gpio_pins_0_13[1].gpio_instance.function_reg ),
    .Y(_181_));
 sky130_fd_sc_hd__nand2b_1 _307_ (.A_N(\gpio_instance_14.enable_reg ),
    .B(\gpio_pins_0_13[0].gpio_instance.function_reg ),
    .Y(_180_));
 sky130_fd_sc_hd__nand2b_1 _308_ (.A_N(\gpio_instance_14.enable_reg ),
    .B(\gpio_instance_15.function_reg ),
    .Y(_179_));
 sky130_fd_sc_hd__nand2b_1 _309_ (.A_N(\gpio_instance_14.enable_reg ),
    .B(\gpio_instance_14.function_reg ),
    .Y(_178_));
 sky130_fd_sc_hd__or2_1 _310_ (.A(\gpio_instance_15.IRQ_INT ),
    .B(\gpio_instance_14.IRQ_INT ),
    .X(net57));
 sky130_fd_sc_hd__o21bai_1 _311_ (.A1(net36),
    .A2(_134_),
    .B1_N(PIN_DATA[14]),
    .Y(_176_));
 sky130_fd_sc_hd__o311a_1 _312_ (.A1(net36),
    .A2(\gpio_instance_14.Data_in ),
    .A3(_134_),
    .B1(_130_),
    .C1(_176_),
    .X(_000_));
 sky130_fd_sc_hd__o211a_1 _313_ (.A1(net36),
    .A2(_134_),
    .B1(_172_),
    .C1(\gpio_instance_14.irq_detected ),
    .X(_001_));
 sky130_fd_sc_hd__o21bai_1 _314_ (.A1(net37),
    .A2(_135_),
    .B1_N(PIN_DATA[15]),
    .Y(_177_));
 sky130_fd_sc_hd__o311a_1 _315_ (.A1(net37),
    .A2(\gpio_instance_15.Data_in ),
    .A3(_135_),
    .B1(_130_),
    .C1(_177_),
    .X(_003_));
 sky130_fd_sc_hd__o211a_1 _316_ (.A1(net37),
    .A2(_135_),
    .B1(_166_),
    .C1(\gpio_instance_15.irq_detected ),
    .X(_004_));
 sky130_fd_sc_hd__inv_2 _317_ (.A(net38),
    .Y(_067_));
 sky130_fd_sc_hd__inv_2 _318_ (.A(net38),
    .Y(_068_));
 sky130_fd_sc_hd__inv_2 _319_ (.A(net38),
    .Y(_069_));
 sky130_fd_sc_hd__inv_2 _320_ (.A(net38),
    .Y(_070_));
 sky130_fd_sc_hd__inv_2 _321_ (.A(net38),
    .Y(_071_));
 sky130_fd_sc_hd__inv_2 _322_ (.A(net38),
    .Y(_072_));
 sky130_fd_sc_hd__inv_2 _323_ (.A(net38),
    .Y(_073_));
 sky130_fd_sc_hd__inv_2 _324_ (.A(net38),
    .Y(_074_));
 sky130_fd_sc_hd__inv_2 _325_ (.A(net38),
    .Y(_075_));
 sky130_fd_sc_hd__inv_2 _326_ (.A(net38),
    .Y(_076_));
 sky130_fd_sc_hd__inv_2 _327_ (.A(net38),
    .Y(_077_));
 sky130_fd_sc_hd__inv_2 _328_ (.A(net38),
    .Y(_078_));
 sky130_fd_sc_hd__inv_2 _329_ (.A(net38),
    .Y(_079_));
 sky130_fd_sc_hd__inv_2 _330_ (.A(net38),
    .Y(_080_));
 sky130_fd_sc_hd__inv_2 _331_ (.A(net38),
    .Y(_081_));
 sky130_fd_sc_hd__inv_2 _332_ (.A(net38),
    .Y(_082_));
 sky130_fd_sc_hd__inv_2 _333_ (.A(net38),
    .Y(_083_));
 sky130_fd_sc_hd__inv_2 _334_ (.A(net38),
    .Y(_084_));
 sky130_fd_sc_hd__inv_2 _335_ (.A(net38),
    .Y(_085_));
 sky130_fd_sc_hd__inv_2 _336_ (.A(net38),
    .Y(_086_));
 sky130_fd_sc_hd__inv_2 _337_ (.A(net38),
    .Y(_087_));
 sky130_fd_sc_hd__inv_2 _338_ (.A(net38),
    .Y(_088_));
 sky130_fd_sc_hd__inv_2 _339_ (.A(net38),
    .Y(_089_));
 sky130_fd_sc_hd__inv_2 _340_ (.A(net38),
    .Y(_090_));
 sky130_fd_sc_hd__inv_2 _341_ (.A(net38),
    .Y(_091_));
 sky130_fd_sc_hd__inv_2 _342_ (.A(net38),
    .Y(_092_));
 sky130_fd_sc_hd__inv_2 _343_ (.A(net38),
    .Y(_093_));
 sky130_fd_sc_hd__inv_2 _344_ (.A(net38),
    .Y(_094_));
 sky130_fd_sc_hd__inv_2 _345_ (.A(net38),
    .Y(_020_));
 sky130_fd_sc_hd__inv_2 _346_ (.A(net38),
    .Y(_021_));
 sky130_fd_sc_hd__inv_2 _347_ (.A(net38),
    .Y(_022_));
 sky130_fd_sc_hd__inv_2 _348_ (.A(net38),
    .Y(_023_));
 sky130_fd_sc_hd__inv_2 _349_ (.A(net38),
    .Y(_024_));
 sky130_fd_sc_hd__inv_2 _350_ (.A(net38),
    .Y(_025_));
 sky130_fd_sc_hd__inv_2 _351_ (.A(net38),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _352_ (.A(net38),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _353_ (.A(net38),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _354_ (.A(net38),
    .Y(_029_));
 sky130_fd_sc_hd__inv_2 _355_ (.A(net38),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _356_ (.A(net38),
    .Y(_031_));
 sky130_fd_sc_hd__inv_2 _357_ (.A(net38),
    .Y(_032_));
 sky130_fd_sc_hd__inv_2 _358_ (.A(net38),
    .Y(_033_));
 sky130_fd_sc_hd__inv_2 _359_ (.A(net38),
    .Y(_034_));
 sky130_fd_sc_hd__inv_2 _360_ (.A(net38),
    .Y(_035_));
 sky130_fd_sc_hd__inv_2 _361_ (.A(net38),
    .Y(_036_));
 sky130_fd_sc_hd__inv_2 _362_ (.A(net38),
    .Y(_037_));
 sky130_fd_sc_hd__inv_2 _363_ (.A(net38),
    .Y(_038_));
 sky130_fd_sc_hd__inv_2 _364_ (.A(net38),
    .Y(_039_));
 sky130_fd_sc_hd__inv_2 _365_ (.A(net38),
    .Y(_040_));
 sky130_fd_sc_hd__inv_2 _366_ (.A(net38),
    .Y(_041_));
 sky130_fd_sc_hd__inv_2 _367_ (.A(net38),
    .Y(_042_));
 sky130_fd_sc_hd__inv_2 _368_ (.A(net38),
    .Y(_043_));
 sky130_fd_sc_hd__inv_2 _369_ (.A(net38),
    .Y(_044_));
 sky130_fd_sc_hd__inv_2 _370_ (.A(net38),
    .Y(_045_));
 sky130_fd_sc_hd__inv_2 _371_ (.A(net38),
    .Y(_046_));
 sky130_fd_sc_hd__inv_2 _372_ (.A(net38),
    .Y(_047_));
 sky130_fd_sc_hd__inv_2 _373_ (.A(net38),
    .Y(_048_));
 sky130_fd_sc_hd__inv_2 _374_ (.A(net38),
    .Y(_049_));
 sky130_fd_sc_hd__inv_2 _375_ (.A(net38),
    .Y(_050_));
 sky130_fd_sc_hd__inv_2 _376_ (.A(net38),
    .Y(_051_));
 sky130_fd_sc_hd__inv_2 _377_ (.A(net38),
    .Y(_052_));
 sky130_fd_sc_hd__inv_2 _378_ (.A(net38),
    .Y(_053_));
 sky130_fd_sc_hd__inv_2 _379_ (.A(net38),
    .Y(_054_));
 sky130_fd_sc_hd__inv_2 _380_ (.A(net38),
    .Y(_055_));
 sky130_fd_sc_hd__inv_2 _381_ (.A(net38),
    .Y(_056_));
 sky130_fd_sc_hd__inv_2 _382_ (.A(net38),
    .Y(_057_));
 sky130_fd_sc_hd__inv_2 _383_ (.A(net38),
    .Y(_058_));
 sky130_fd_sc_hd__inv_2 _384_ (.A(net38),
    .Y(_059_));
 sky130_fd_sc_hd__inv_2 _385_ (.A(net38),
    .Y(_060_));
 sky130_fd_sc_hd__inv_2 _386_ (.A(net38),
    .Y(_061_));
 sky130_fd_sc_hd__inv_2 _387_ (.A(net38),
    .Y(_062_));
 sky130_fd_sc_hd__inv_2 _388_ (.A(net38),
    .Y(_063_));
 sky130_fd_sc_hd__inv_2 _389_ (.A(net38),
    .Y(_064_));
 sky130_fd_sc_hd__inv_2 _390_ (.A(net38),
    .Y(_065_));
 sky130_fd_sc_hd__dfrtp_1 _391_ (.CLK(clknet_3_1__leaf_clk),
    .D(_119_),
    .RESET_B(_066_),
    .Q(\gpio_instance_14.PIN_DATA_prev ));
 sky130_fd_sc_hd__dfrtp_4 _392_ (.CLK(clknet_3_6__leaf_clk),
    .D(net17),
    .RESET_B(_067_),
    .Q(\gpio_instance_14.enable_reg ));
 sky130_fd_sc_hd__dfrtp_1 _393_ (.CLK(clknet_3_1__leaf_clk),
    .D(_001_),
    .RESET_B(_068_),
    .Q(\gpio_instance_14.IRQ_INT ));
 sky130_fd_sc_hd__dfrtp_1 _394_ (.CLK(clknet_3_0__leaf_clk),
    .D(_002_),
    .RESET_B(_069_),
    .Q(\gpio_instance_14.Pin_out ));
 sky130_fd_sc_hd__dfrtp_1 _395_ (.CLK(clknet_3_0__leaf_clk),
    .D(\gpio_instance_14.Function ),
    .RESET_B(_070_),
    .Q(\gpio_instance_14.function_reg ));
 sky130_fd_sc_hd__dfrtp_1 _396_ (.CLK(clknet_3_0__leaf_clk),
    .D(_000_),
    .RESET_B(_071_),
    .Q(\gpio_instance_14.Data_in ));
 sky130_fd_sc_hd__dfrtp_1 _397_ (.CLK(clknet_3_0__leaf_clk),
    .D(net36),
    .RESET_B(_072_),
    .Q(\gpio_instance_14.pin_change_mask_reg ));
 sky130_fd_sc_hd__dfrtp_1 _398_ (.CLK(clknet_3_1__leaf_clk),
    .D(_120_),
    .RESET_B(_073_),
    .Q(\gpio_instance_14.irq_detected ));
 sky130_fd_sc_hd__dfrtp_1 _399_ (.CLK(clknet_3_1__leaf_clk),
    .D(net34),
    .RESET_B(_074_),
    .Q(\gpio_instance_14.int_mask_reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _400_ (.CLK(clknet_3_1__leaf_clk),
    .D(net35),
    .RESET_B(_075_),
    .Q(\gpio_instance_14.int_mask_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _401_ (.CLK(clknet_3_1__leaf_clk),
    .D(_121_),
    .RESET_B(_076_),
    .Q(\gpio_instance_15.PIN_DATA_prev ));
 sky130_fd_sc_hd__dfrtp_1 _402_ (.CLK(clknet_3_1__leaf_clk),
    .D(_004_),
    .RESET_B(_077_),
    .Q(\gpio_instance_15.IRQ_INT ));
 sky130_fd_sc_hd__dfrtp_1 _403_ (.CLK(clknet_3_4__leaf_clk),
    .D(_005_),
    .RESET_B(_078_),
    .Q(\gpio_instance_15.Pin_out ));
 sky130_fd_sc_hd__dfrtp_1 _404_ (.CLK(clknet_3_4__leaf_clk),
    .D(\gpio_instance_15.Function ),
    .RESET_B(_079_),
    .Q(\gpio_instance_15.function_reg ));
 sky130_fd_sc_hd__dfrtp_1 _405_ (.CLK(clknet_3_4__leaf_clk),
    .D(_003_),
    .RESET_B(_080_),
    .Q(\gpio_instance_15.Data_in ));
 sky130_fd_sc_hd__dfrtp_1 _406_ (.CLK(clknet_3_0__leaf_clk),
    .D(_122_),
    .RESET_B(_081_),
    .Q(\gpio_instance_14.pin_value ));
 sky130_fd_sc_hd__dfrtp_1 _407_ (.CLK(clknet_3_4__leaf_clk),
    .D(net37),
    .RESET_B(_082_),
    .Q(\gpio_instance_15.pin_change_mask_reg ));
 sky130_fd_sc_hd__dfrtp_1 _408_ (.CLK(clknet_3_1__leaf_clk),
    .D(_123_),
    .RESET_B(_083_),
    .Q(\gpio_instance_15.irq_detected ));
 sky130_fd_sc_hd__dfrtp_1 _409_ (.CLK(clknet_3_0__leaf_clk),
    .D(_124_),
    .RESET_B(_084_),
    .Q(\gpio_pins_0_13[9].gpio_instance.pin_value ));
 sky130_fd_sc_hd__dfrtp_1 _410_ (.CLK(clknet_3_5__leaf_clk),
    .D(_006_),
    .RESET_B(_085_),
    .Q(\gpio_pins_0_13[0].gpio_instance.Pin_out ));
 sky130_fd_sc_hd__dfrtp_1 _411_ (.CLK(clknet_3_5__leaf_clk),
    .D(net18),
    .RESET_B(_086_),
    .Q(\gpio_pins_0_13[0].gpio_instance.function_reg ));
 sky130_fd_sc_hd__dfrtp_1 _412_ (.CLK(clknet_3_4__leaf_clk),
    .D(_125_),
    .RESET_B(_087_),
    .Q(\gpio_instance_15.pin_value ));
 sky130_fd_sc_hd__dfrtp_1 _413_ (.CLK(clknet_3_2__leaf_clk),
    .D(_011_),
    .RESET_B(_088_),
    .Q(\gpio_pins_0_13[1].gpio_instance.Pin_out ));
 sky130_fd_sc_hd__dfrtp_1 _414_ (.CLK(clknet_3_2__leaf_clk),
    .D(net25),
    .RESET_B(_089_),
    .Q(\gpio_pins_0_13[1].gpio_instance.function_reg ));
 sky130_fd_sc_hd__dfrtp_1 _415_ (.CLK(clknet_3_3__leaf_clk),
    .D(_126_),
    .RESET_B(_090_),
    .Q(\gpio_pins_0_13[13].gpio_instance.Data_in ));
 sky130_fd_sc_hd__dfrtp_1 _416_ (.CLK(clknet_3_3__leaf_clk),
    .D(_127_),
    .RESET_B(_091_),
    .Q(\gpio_pins_0_13[13].gpio_instance.pin_value ));
 sky130_fd_sc_hd__dfrtp_1 _417_ (.CLK(clknet_3_3__leaf_clk),
    .D(_012_),
    .RESET_B(_092_),
    .Q(\gpio_pins_0_13[2].gpio_instance.Pin_out ));
 sky130_fd_sc_hd__dfrtp_1 _418_ (.CLK(clknet_3_6__leaf_clk),
    .D(net26),
    .RESET_B(_093_),
    .Q(\gpio_pins_0_13[2].gpio_instance.function_reg ));
 sky130_fd_sc_hd__dfrtp_1 _419_ (.CLK(clknet_3_2__leaf_clk),
    .D(_128_),
    .RESET_B(_094_),
    .Q(\gpio_pins_0_13[1].gpio_instance.Data_in ));
 sky130_fd_sc_hd__dfrtp_1 _420_ (.CLK(clknet_3_2__leaf_clk),
    .D(_095_),
    .RESET_B(_020_),
    .Q(\gpio_pins_0_13[1].gpio_instance.pin_value ));
 sky130_fd_sc_hd__dfrtp_1 _421_ (.CLK(clknet_3_4__leaf_clk),
    .D(_013_),
    .RESET_B(_021_),
    .Q(\gpio_pins_0_13[3].gpio_instance.Pin_out ));
 sky130_fd_sc_hd__dfrtp_1 _422_ (.CLK(clknet_3_4__leaf_clk),
    .D(net27),
    .RESET_B(_022_),
    .Q(\gpio_pins_0_13[3].gpio_instance.function_reg ));
 sky130_fd_sc_hd__dfrtp_1 _423_ (.CLK(clknet_3_6__leaf_clk),
    .D(_096_),
    .RESET_B(_023_),
    .Q(\gpio_pins_0_13[2].gpio_instance.Data_in ));
 sky130_fd_sc_hd__dfrtp_1 _424_ (.CLK(clknet_3_3__leaf_clk),
    .D(_097_),
    .RESET_B(_024_),
    .Q(\gpio_pins_0_13[2].gpio_instance.pin_value ));
 sky130_fd_sc_hd__dfrtp_1 _425_ (.CLK(clknet_3_7__leaf_clk),
    .D(_014_),
    .RESET_B(_025_),
    .Q(\gpio_pins_0_13[4].gpio_instance.Pin_out ));
 sky130_fd_sc_hd__dfrtp_1 _426_ (.CLK(clknet_3_7__leaf_clk),
    .D(net28),
    .RESET_B(_026_),
    .Q(\gpio_pins_0_13[4].gpio_instance.function_reg ));
 sky130_fd_sc_hd__dfrtp_1 _427_ (.CLK(clknet_3_5__leaf_clk),
    .D(_098_),
    .RESET_B(_027_),
    .Q(\gpio_pins_0_13[3].gpio_instance.Data_in ));
 sky130_fd_sc_hd__dfrtp_1 _428_ (.CLK(clknet_3_5__leaf_clk),
    .D(_099_),
    .RESET_B(_028_),
    .Q(\gpio_pins_0_13[3].gpio_instance.pin_value ));
 sky130_fd_sc_hd__dfrtp_1 _429_ (.CLK(clknet_3_0__leaf_clk),
    .D(_015_),
    .RESET_B(_029_),
    .Q(\gpio_pins_0_13[5].gpio_instance.Pin_out ));
 sky130_fd_sc_hd__dfrtp_1 _430_ (.CLK(clknet_3_0__leaf_clk),
    .D(net29),
    .RESET_B(_030_),
    .Q(\gpio_pins_0_13[5].gpio_instance.function_reg ));
 sky130_fd_sc_hd__dfrtp_1 _431_ (.CLK(clknet_3_7__leaf_clk),
    .D(_100_),
    .RESET_B(_031_),
    .Q(\gpio_pins_0_13[4].gpio_instance.Data_in ));
 sky130_fd_sc_hd__dfrtp_1 _432_ (.CLK(clknet_3_6__leaf_clk),
    .D(_101_),
    .RESET_B(_032_),
    .Q(\gpio_pins_0_13[4].gpio_instance.pin_value ));
 sky130_fd_sc_hd__dfrtp_1 _433_ (.CLK(clknet_3_5__leaf_clk),
    .D(_016_),
    .RESET_B(_033_),
    .Q(\gpio_pins_0_13[6].gpio_instance.Pin_out ));
 sky130_fd_sc_hd__dfrtp_1 _434_ (.CLK(clknet_3_5__leaf_clk),
    .D(net30),
    .RESET_B(_034_),
    .Q(\gpio_pins_0_13[6].gpio_instance.function_reg ));
 sky130_fd_sc_hd__dfrtp_1 _435_ (.CLK(clknet_3_3__leaf_clk),
    .D(_102_),
    .RESET_B(_035_),
    .Q(\gpio_pins_0_13[5].gpio_instance.Data_in ));
 sky130_fd_sc_hd__dfrtp_1 _436_ (.CLK(clknet_3_0__leaf_clk),
    .D(_103_),
    .RESET_B(_036_),
    .Q(\gpio_pins_0_13[5].gpio_instance.pin_value ));
 sky130_fd_sc_hd__dfrtp_1 _437_ (.CLK(clknet_3_6__leaf_clk),
    .D(_017_),
    .RESET_B(_037_),
    .Q(\gpio_pins_0_13[7].gpio_instance.Pin_out ));
 sky130_fd_sc_hd__dfrtp_1 _438_ (.CLK(clknet_3_6__leaf_clk),
    .D(net31),
    .RESET_B(_038_),
    .Q(\gpio_pins_0_13[7].gpio_instance.function_reg ));
 sky130_fd_sc_hd__dfrtp_1 _439_ (.CLK(clknet_3_5__leaf_clk),
    .D(_104_),
    .RESET_B(_039_),
    .Q(\gpio_pins_0_13[6].gpio_instance.Data_in ));
 sky130_fd_sc_hd__dfrtp_1 _440_ (.CLK(clknet_3_5__leaf_clk),
    .D(_105_),
    .RESET_B(_040_),
    .Q(\gpio_pins_0_13[6].gpio_instance.pin_value ));
 sky130_fd_sc_hd__dfrtp_1 _441_ (.CLK(clknet_3_7__leaf_clk),
    .D(_018_),
    .RESET_B(_041_),
    .Q(\gpio_pins_0_13[8].gpio_instance.Pin_out ));
 sky130_fd_sc_hd__dfrtp_1 _442_ (.CLK(clknet_3_7__leaf_clk),
    .D(net32),
    .RESET_B(_042_),
    .Q(\gpio_pins_0_13[8].gpio_instance.function_reg ));
 sky130_fd_sc_hd__dfrtp_1 _443_ (.CLK(clknet_3_6__leaf_clk),
    .D(_106_),
    .RESET_B(_043_),
    .Q(\gpio_pins_0_13[7].gpio_instance.Data_in ));
 sky130_fd_sc_hd__dfrtp_1 _444_ (.CLK(clknet_3_6__leaf_clk),
    .D(_107_),
    .RESET_B(_044_),
    .Q(\gpio_pins_0_13[7].gpio_instance.pin_value ));
 sky130_fd_sc_hd__dfrtp_1 _445_ (.CLK(clknet_3_0__leaf_clk),
    .D(_108_),
    .RESET_B(_045_),
    .Q(\gpio_pins_0_13[9].gpio_instance.Data_in ));
 sky130_fd_sc_hd__dfrtp_1 _446_ (.CLK(clknet_3_0__leaf_clk),
    .D(_019_),
    .RESET_B(_046_),
    .Q(\gpio_pins_0_13[9].gpio_instance.Pin_out ));
 sky130_fd_sc_hd__dfrtp_1 _447_ (.CLK(clknet_3_0__leaf_clk),
    .D(net33),
    .RESET_B(_047_),
    .Q(\gpio_pins_0_13[9].gpio_instance.function_reg ));
 sky130_fd_sc_hd__dfrtp_1 _448_ (.CLK(clknet_3_7__leaf_clk),
    .D(_109_),
    .RESET_B(_048_),
    .Q(\gpio_pins_0_13[8].gpio_instance.Data_in ));
 sky130_fd_sc_hd__dfrtp_1 _449_ (.CLK(clknet_3_7__leaf_clk),
    .D(_110_),
    .RESET_B(_049_),
    .Q(\gpio_pins_0_13[8].gpio_instance.pin_value ));
 sky130_fd_sc_hd__dfrtp_1 _450_ (.CLK(clknet_3_3__leaf_clk),
    .D(_007_),
    .RESET_B(_050_),
    .Q(\gpio_pins_0_13[10].gpio_instance.Pin_out ));
 sky130_fd_sc_hd__dfrtp_1 _451_ (.CLK(clknet_3_2__leaf_clk),
    .D(net19),
    .RESET_B(_051_),
    .Q(\gpio_pins_0_13[10].gpio_instance.function_reg ));
 sky130_fd_sc_hd__dfrtp_1 _452_ (.CLK(clknet_3_5__leaf_clk),
    .D(_111_),
    .RESET_B(_052_),
    .Q(\gpio_pins_0_13[0].gpio_instance.Data_in ));
 sky130_fd_sc_hd__dfrtp_1 _453_ (.CLK(clknet_3_5__leaf_clk),
    .D(_112_),
    .RESET_B(_053_),
    .Q(\gpio_pins_0_13[0].gpio_instance.pin_value ));
 sky130_fd_sc_hd__dfrtp_1 _454_ (.CLK(clknet_3_2__leaf_clk),
    .D(_008_),
    .RESET_B(_054_),
    .Q(\gpio_pins_0_13[11].gpio_instance.Pin_out ));
 sky130_fd_sc_hd__dfrtp_1 _455_ (.CLK(clknet_3_2__leaf_clk),
    .D(net20),
    .RESET_B(_055_),
    .Q(\gpio_pins_0_13[11].gpio_instance.function_reg ));
 sky130_fd_sc_hd__dfrtp_1 _456_ (.CLK(clknet_3_2__leaf_clk),
    .D(_113_),
    .RESET_B(_056_),
    .Q(\gpio_pins_0_13[10].gpio_instance.Data_in ));
 sky130_fd_sc_hd__dfrtp_1 _457_ (.CLK(clknet_3_3__leaf_clk),
    .D(_114_),
    .RESET_B(_057_),
    .Q(\gpio_pins_0_13[10].gpio_instance.pin_value ));
 sky130_fd_sc_hd__dfrtp_1 _458_ (.CLK(clknet_3_7__leaf_clk),
    .D(_009_),
    .RESET_B(_058_),
    .Q(\gpio_pins_0_13[12].gpio_instance.Pin_out ));
 sky130_fd_sc_hd__dfrtp_1 _459_ (.CLK(clknet_3_7__leaf_clk),
    .D(net21),
    .RESET_B(_059_),
    .Q(\gpio_pins_0_13[12].gpio_instance.function_reg ));
 sky130_fd_sc_hd__dfrtp_1 _460_ (.CLK(clknet_3_2__leaf_clk),
    .D(_115_),
    .RESET_B(_060_),
    .Q(\gpio_pins_0_13[11].gpio_instance.Data_in ));
 sky130_fd_sc_hd__dfrtp_1 _461_ (.CLK(clknet_3_2__leaf_clk),
    .D(_116_),
    .RESET_B(_061_),
    .Q(\gpio_pins_0_13[11].gpio_instance.pin_value ));
 sky130_fd_sc_hd__dfrtp_1 _462_ (.CLK(clknet_3_2__leaf_clk),
    .D(_010_),
    .RESET_B(_062_),
    .Q(\gpio_pins_0_13[13].gpio_instance.Pin_out ));
 sky130_fd_sc_hd__dfrtp_1 _463_ (.CLK(clknet_3_3__leaf_clk),
    .D(net22),
    .RESET_B(_063_),
    .Q(\gpio_pins_0_13[13].gpio_instance.function_reg ));
 sky130_fd_sc_hd__dfrtp_1 _464_ (.CLK(clknet_3_7__leaf_clk),
    .D(_117_),
    .RESET_B(_064_),
    .Q(\gpio_pins_0_13[12].gpio_instance.Data_in ));
 sky130_fd_sc_hd__dfrtp_1 _465_ (.CLK(clknet_3_7__leaf_clk),
    .D(_118_),
    .RESET_B(_065_),
    .Q(\gpio_pins_0_13[12].gpio_instance.pin_value ));
 sky130_fd_sc_hd__clkbuf_1 _466_ (.A(\gpio_pins_0_13[0].gpio_instance.Data_in ),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 _467_ (.A(\gpio_pins_0_13[1].gpio_instance.Data_in ),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 _468_ (.A(\gpio_pins_0_13[2].gpio_instance.Data_in ),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 _469_ (.A(\gpio_pins_0_13[3].gpio_instance.Data_in ),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 _470_ (.A(\gpio_pins_0_13[4].gpio_instance.Data_in ),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 _471_ (.A(\gpio_pins_0_13[5].gpio_instance.Data_in ),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 _472_ (.A(\gpio_pins_0_13[6].gpio_instance.Data_in ),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 _473_ (.A(\gpio_pins_0_13[7].gpio_instance.Data_in ),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 _474_ (.A(\gpio_pins_0_13[8].gpio_instance.Data_in ),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 _475_ (.A(\gpio_pins_0_13[9].gpio_instance.Data_in ),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 _476_ (.A(\gpio_pins_0_13[10].gpio_instance.Data_in ),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 _477_ (.A(\gpio_pins_0_13[11].gpio_instance.Data_in ),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 _478_ (.A(\gpio_pins_0_13[12].gpio_instance.Data_in ),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 _479_ (.A(\gpio_pins_0_13[13].gpio_instance.Data_in ),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 _480_ (.A(\gpio_instance_14.Data_in ),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 _481_ (.A(\gpio_instance_15.Data_in ),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 _482_ (.A(\gpio_instance_14.IRQ_INT ),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 _483_ (.A(\gpio_instance_15.IRQ_INT ),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 _484_ (.A(\gpio_pins_0_13[0].gpio_instance.Pin_out ),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 _485_ (.A(\gpio_pins_0_13[1].gpio_instance.Pin_out ),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 _486_ (.A(\gpio_pins_0_13[2].gpio_instance.Pin_out ),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 _487_ (.A(\gpio_pins_0_13[3].gpio_instance.Pin_out ),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 _488_ (.A(\gpio_pins_0_13[4].gpio_instance.Pin_out ),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 _489_ (.A(\gpio_pins_0_13[5].gpio_instance.Pin_out ),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 _490_ (.A(\gpio_pins_0_13[6].gpio_instance.Pin_out ),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 _491_ (.A(\gpio_pins_0_13[7].gpio_instance.Pin_out ),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 _492_ (.A(\gpio_pins_0_13[8].gpio_instance.Pin_out ),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 _493_ (.A(\gpio_pins_0_13[9].gpio_instance.Pin_out ),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 _494_ (.A(\gpio_pins_0_13[10].gpio_instance.Pin_out ),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 _495_ (.A(\gpio_pins_0_13[11].gpio_instance.Pin_out ),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 _496_ (.A(\gpio_pins_0_13[12].gpio_instance.Pin_out ),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 _497_ (.A(\gpio_pins_0_13[13].gpio_instance.Pin_out ),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 _498_ (.A(\gpio_instance_14.Pin_out ),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 _499_ (.A(\gpio_instance_15.Pin_out ),
    .X(net64));
 sky130_fd_sc_hd__ebufn_2 _500_ (.A(\gpio_instance_14.pin_value ),
    .TE_B(_178_),
    .Z(PIN_DATA[14]));
 sky130_fd_sc_hd__ebufn_2 _501_ (.A(\gpio_instance_15.pin_value ),
    .TE_B(_179_),
    .Z(PIN_DATA[15]));
 sky130_fd_sc_hd__ebufn_1 _502_ (.A(\gpio_pins_0_13[0].gpio_instance.pin_value ),
    .TE_B(_180_),
    .Z(PIN_DATA[0]));
 sky130_fd_sc_hd__ebufn_1 _503_ (.A(\gpio_pins_0_13[1].gpio_instance.pin_value ),
    .TE_B(_181_),
    .Z(PIN_DATA[1]));
 sky130_fd_sc_hd__ebufn_1 _504_ (.A(\gpio_pins_0_13[2].gpio_instance.pin_value ),
    .TE_B(_182_),
    .Z(PIN_DATA[2]));
 sky130_fd_sc_hd__ebufn_1 _505_ (.A(\gpio_pins_0_13[3].gpio_instance.pin_value ),
    .TE_B(_183_),
    .Z(PIN_DATA[3]));
 sky130_fd_sc_hd__ebufn_1 _506_ (.A(\gpio_pins_0_13[4].gpio_instance.pin_value ),
    .TE_B(_184_),
    .Z(PIN_DATA[4]));
 sky130_fd_sc_hd__ebufn_1 _507_ (.A(\gpio_pins_0_13[5].gpio_instance.pin_value ),
    .TE_B(_185_),
    .Z(PIN_DATA[5]));
 sky130_fd_sc_hd__ebufn_1 _508_ (.A(\gpio_pins_0_13[6].gpio_instance.pin_value ),
    .TE_B(_186_),
    .Z(PIN_DATA[6]));
 sky130_fd_sc_hd__ebufn_1 _509_ (.A(\gpio_pins_0_13[7].gpio_instance.pin_value ),
    .TE_B(_187_),
    .Z(PIN_DATA[7]));
 sky130_fd_sc_hd__ebufn_1 _510_ (.A(\gpio_pins_0_13[8].gpio_instance.pin_value ),
    .TE_B(_188_),
    .Z(PIN_DATA[8]));
 sky130_fd_sc_hd__ebufn_1 _511_ (.A(\gpio_pins_0_13[9].gpio_instance.pin_value ),
    .TE_B(_189_),
    .Z(PIN_DATA[9]));
 sky130_fd_sc_hd__ebufn_1 _512_ (.A(\gpio_pins_0_13[10].gpio_instance.pin_value ),
    .TE_B(_190_),
    .Z(PIN_DATA[10]));
 sky130_fd_sc_hd__ebufn_1 _513_ (.A(\gpio_pins_0_13[11].gpio_instance.pin_value ),
    .TE_B(_191_),
    .Z(PIN_DATA[11]));
 sky130_fd_sc_hd__ebufn_1 _514_ (.A(\gpio_pins_0_13[12].gpio_instance.pin_value ),
    .TE_B(_192_),
    .Z(PIN_DATA[12]));
 sky130_fd_sc_hd__ebufn_1 _515_ (.A(\gpio_pins_0_13[13].gpio_instance.pin_value ),
    .TE_B(_193_),
    .Z(PIN_DATA[13]));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_170 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(Data_out[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(Data_out[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(Data_out[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(Data_out[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(Data_out[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(Data_out[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(Data_out[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(Data_out[1]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(Data_out[2]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(Data_out[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(Data_out[4]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(Data_out[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(Data_out[6]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(Data_out[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(Data_out[8]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(Data_out[9]),
    .X(net16));
 sky130_fd_sc_hd__buf_8 input17 (.A(Enable),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(Function[0]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(Function[10]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(Function[11]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(Function[12]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(Function[13]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(Function[14]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(Function[15]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(Function[1]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(Function[2]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(Function[3]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(Function[4]),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 input29 (.A(Function[5]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input30 (.A(Function[6]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(Function[7]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(Function[8]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(Function[9]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(Int_Mask[0]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(Int_Mask[1]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(Pin_Change_Mask[14]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(Pin_Change_Mask[15]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_16 input38 (.A(reset),
    .X(net38));
 sky130_fd_sc_hd__buf_1 output39 (.A(net39),
    .X(Data_in[0]));
 sky130_fd_sc_hd__buf_1 output40 (.A(net40),
    .X(Data_in[10]));
 sky130_fd_sc_hd__buf_1 output41 (.A(net41),
    .X(Data_in[11]));
 sky130_fd_sc_hd__buf_1 output42 (.A(net42),
    .X(Data_in[12]));
 sky130_fd_sc_hd__buf_1 output43 (.A(net43),
    .X(Data_in[13]));
 sky130_fd_sc_hd__buf_1 output44 (.A(net44),
    .X(Data_in[14]));
 sky130_fd_sc_hd__buf_1 output45 (.A(net45),
    .X(Data_in[15]));
 sky130_fd_sc_hd__buf_1 output46 (.A(net46),
    .X(Data_in[1]));
 sky130_fd_sc_hd__buf_1 output47 (.A(net47),
    .X(Data_in[2]));
 sky130_fd_sc_hd__buf_1 output48 (.A(net48),
    .X(Data_in[3]));
 sky130_fd_sc_hd__buf_1 output49 (.A(net49),
    .X(Data_in[4]));
 sky130_fd_sc_hd__buf_1 output50 (.A(net50),
    .X(Data_in[5]));
 sky130_fd_sc_hd__buf_1 output51 (.A(net51),
    .X(Data_in[6]));
 sky130_fd_sc_hd__buf_1 output52 (.A(net52),
    .X(Data_in[7]));
 sky130_fd_sc_hd__buf_1 output53 (.A(net53),
    .X(Data_in[8]));
 sky130_fd_sc_hd__buf_1 output54 (.A(net54),
    .X(Data_in[9]));
 sky130_fd_sc_hd__buf_1 output55 (.A(net55),
    .X(IRQ_INT[0]));
 sky130_fd_sc_hd__buf_1 output56 (.A(net56),
    .X(IRQ_INT[1]));
 sky130_fd_sc_hd__buf_1 output57 (.A(net57),
    .X(IRQ_PIN_CHANGE));
 sky130_fd_sc_hd__buf_1 output58 (.A(net58),
    .X(Pin_out[0]));
 sky130_fd_sc_hd__buf_1 output59 (.A(net59),
    .X(Pin_out[10]));
 sky130_fd_sc_hd__buf_1 output60 (.A(net60),
    .X(Pin_out[11]));
 sky130_fd_sc_hd__buf_1 output61 (.A(net61),
    .X(Pin_out[12]));
 sky130_fd_sc_hd__buf_1 output62 (.A(net62),
    .X(Pin_out[13]));
 sky130_fd_sc_hd__buf_1 output63 (.A(net63),
    .X(Pin_out[14]));
 sky130_fd_sc_hd__buf_1 output64 (.A(net64),
    .X(Pin_out[15]));
 sky130_fd_sc_hd__buf_1 output65 (.A(net65),
    .X(Pin_out[1]));
 sky130_fd_sc_hd__buf_1 output66 (.A(net66),
    .X(Pin_out[2]));
 sky130_fd_sc_hd__buf_1 output67 (.A(net67),
    .X(Pin_out[3]));
 sky130_fd_sc_hd__buf_1 output68 (.A(net68),
    .X(Pin_out[4]));
 sky130_fd_sc_hd__buf_1 output69 (.A(net69),
    .X(Pin_out[5]));
 sky130_fd_sc_hd__buf_1 output70 (.A(net70),
    .X(Pin_out[6]));
 sky130_fd_sc_hd__buf_1 output71 (.A(net71),
    .X(Pin_out[7]));
 sky130_fd_sc_hd__buf_1 output72 (.A(net72),
    .X(Pin_out[8]));
 sky130_fd_sc_hd__buf_1 output73 (.A(net73),
    .X(Pin_out[9]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__bufinv_16 clkload0 (.A(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload1 (.A(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__bufinv_16 clkload2 (.A(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload3 (.A(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload4 (.A(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__bufinv_16 clkload5 (.A(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload6 (.A(clknet_3_7__leaf_clk));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_191 ();
endmodule
